PK   [�T;m7�  ��     cirkitFile.json�]K��6�+[�UT/��fU>d�Z��ϔ���*�4KIv�.��H����t��C|�-��h _?� ȯ�<��m��]��?g�~��N��N��<��\?����v~��ɓ����W�;8����ݧ��6��I�Jy����X W���(X�e��4[0�����Ǯ��KX�_�$�i��T&��Xe���Bi�|�4}u�Ӳ���mˈ�#8�.1-���n�"\u��7l�#L�N�W����>%��V(�樶�m���#QmK�)����"�E 3��`YG�\�%SJĚ1��(�`�0r��g @M�|	3>�e1����b)u��|�_E�����"-��~�f�{��i\���.-_�,N�E�Wփ�<0�*�I�8��\p�5_� jTܐ��!@n\�^�ƭa��U��6ʒ2M�H�@��(�#�\��L���H��L��8�Ƙ�Q�-|-˒�J��M�֪��V����d�e�ą��g�@M��z�]	d}d�$��\���	��B��8�>����W�>�q�����c��*�+~���i�����uTݯ* ��uH��C��@��0��&��1M�����-�>��{���uH�� Y��d� ��PU�	)`4̤{1زӴ7�e�$Yi�'�T �{�:$y�� ��0��}(�t�"�o�4�5���[�AM�0��}����ĸ��>��e_��aD��3��FJ1-��Ġ��1��_E��T|���`��`�v�V_�6���>�n�
�L��qq<�?qA�"J.��"I�(�E$\t9�n�\�,1	Ұa$#�8A�FҌ���&�13���0C�)s̉l0�悦S�d�����FM3Ćf�c��4(�& 
%[,h�	AN��B�b�.�AC����!��"�+7tC��|B�v�e�Н�.�.èn�pFpCg u�����Y�eu�M��	�{!�2쯁;1\Q�[d��$�"pǃ`\�=5p�c�b¶A� <,lS����¶9�<,l�b���6��aa[�\�;��<��>4�Ь?�|��\�@���\�i}.�j�.���!9d�d�6;�d�L��p.���$�H�D$\4	C�%�Axi��h��h��h �h�h �h0�h@�hP�iP̉l0�9�9�9�9�9�9�9���Q(A�bA�bA�bA�bA�bA�b1�bp��e��d;�� ���v<�A����x.��'���@��x.è�&��\�QM����l�sF4��o2��v<�aM��{kh��e�WC��x.Þ�l���d;�����x. L�� <,0َ���d{/p��eu�d;�� ���v<�Aԁ��\��v<���6����P�k����&�L'_�y���l�e�����.O�|��u�q=MQWM1a��ۡ���f�v�5v�jմD-�PM3Tt�kա2���Q���}McT��4f��;�wz�N���׶�ܤm�ۀ��t�ڛ������e�d��oJ���{�o�9�������>j�4F��ל�y�^�����8p��9��iw9�^-�������� ��F�0c�F^���;���t�6�٧��,�'۴+���
y��Ók'2A 2A 2'A 25A 2CA 2Q�/�-�x	�i�^	n���K�Mb�%��2�Ni���l��Mp" �ǄN�L?bE@�$��@�t��~*��H�)̨��M_w�b����D�f��.f�&��.^��zE�Iz/6K��H����AxP �ېI�E��@2�H.�@�հ(D�/"P��DZ�L���x`���00�n��!�I�/6獅!:�M���p��$O��������n�*�����u�������-v�S�s�F���,]d�f������u{�1��A�#��Q:ЋL����Rm8��L-r��Em~���6��5���<�0�ï�!&�±�w@�I�6�(�mQ��(�\��GM@�!Fŋ��~�����X��0%�!��2�Zy��S6PXll"z,5��?�>C��!�F?�΁����:��?̪�/�c������Ы���}`�^���� �5�`�0���;�����Vؠ��}�z�S�l�[���`�Ћ�v��z��]_<�ڏ�>G��﵌������nxyS�l�����t`ߚ�`�3������u��[���������m�@����(y2����0:=���~L��o�7��c��W��"w���f��l��w�|Ȣ�}<�i�SQ��t9|:P9��u�p�0�2���sѿ�pQq֋�ŉd�j糋#/�Y���w5����)�b�C����(�GWC�����(�p��a�t� ��ě�%X+03���Y&�^���,K�n������d���>%�~E;��}��hK��.*��\�'��}c�~�N`�����u�H�K��N#��!��Y����>in��v��-�m^���Ҡߘ�^1�>�Y��N%������s�o~ҝw �x�r���B����!�:u{A�{ú����67���%���Q�.����m�,����Z�V���q�5JXU��E�*��"Q�v���d�HUE�]UEQ�HWE�]WEq������}f�>�;�N�f�6U�iW;k�;�k	;	k�	;u��{�N�U.ד�f�ȳ$]��]�_����࠹dv�VL�U���� YiH���@e�._=�)?f�1�d�C�>�f�t���=9������|���u��<�����m-A�u4����GN�13�/OLdY;Mx���-��d$��ʲ@.,H�2��U(ujVZ������l�eP~b:��k+{R�69��G�u��dUo>L��E0�GO�
���Dj_I䭣�ub_��p�m�-u��O'<��>y�]��{�M�1 ��xxU<�����=���ġ�D��:�7:⣓|�塴�L��3�f8��t�}%��oI�+q��)��:�i�&���Y΀t<�c-�Hw��ڙ�z���iG��tm~qg�m~�t-~�`��u�=6�����ᘮw?g��4�l�f�m.c��e��q>�R��z��5�����J������~�Yt~��][�4���?�����e:yX%�}f�Y��z�^l��<��q�g�]�ó^�S�=���ᘻ7��[�&����4Y����/���ձ=�K�p�B���\rV�o43ٸ0:M����B.�8�"
�q����$lT�8Z�(^4}'(����E�����iЀ� O�Ъz8���g�R&�L#?uMV�hkU�LO#632���ӓ���zf�
cc���.��y��Q�gvib�S��Ƨ,��C+��!+��4�fƤ��͹%e��jZb�#TrƸ6��uP��+��)u����=���ԁ)����nh��pxƜ"�aS���6U�`�EXjԩ�jiT�Pv,O
U��^��Q�J�N~��^� ��R�X[�=�V�G��:U�w��U���!W�L��U��"�nfS���/�j$Y#ʖS�U��K,REՅn!�fYŪ�|<�Rsy6)*�FE�Z�~��{\9â*�W�*2�J��R3)bf#�@j^zEi�:����M혔�����h��bd.:�I��
2˾��O� u8Q����UDT��g��z���ń:)G��y�E'M�z�K-K�����5��(���-Z��K���R1*m��JA*�R�Дzb*Bs��j����4)2������ܵ�^�-u�05��F�vIg�\e��5F����
M`�,�I��D1a��K��e�hbt��j��e��7�,FWMj��|��O����s�dv),��+������������)`�(��e^�����L6�.7{��TZ�eT�J���]efӅE��XKťu���B�`i�8aL�T�Mp�N� ���*�F�N����	��GC�py��q�X8��M�B��Bc͟m�����:��h�^8���C�{ƫg�Y!���X�Ɗ3d�5k�^g��%��,���Z�g���?��/�q��u)������:�����wN��d�h������(z����[�M{y�N8����R�,�Љ��[o��s��������e��z�
>��wO>���
�:s1�6�ꧣ�v�qYm�%;��ĉ����䛅T�UQN�C�I�C��:thBG��]��+���JV[����:5:"Rt�W�C� t4�j�ҫi��T�d����3�wC��n�vO;�m؀�8o��nx�R��C����-5<�x���G��Q�wL����A���C���u��P���I&��^�]��F��/�t� <$):^xD0�� ��>�G:��n��َ��I6c��l�Q@'>�dm��,�`����<�p�F�]�w{�B�L����V��[��7*B:x�!)<^Th<�d�-�6B�d�=�~�Ao=�F�T�nCã
�x��u2�	���r���f�@7ڨ��v��T�!2�Y�l�Z��z�A�	�g@n	R�cD>,2U�G��T�	�1dWmn`h:n:���MG�7 �����F���m��Fn@2*�d7�lGv��F���R8,�������!�1dw43���j|pZ3c^�B13M�������d�t��6�$[���n�5�?1����ҍ�h�Ͷz2�ʣ����3ӣ���D�7.P�*R��n�ͤ�I�m3�����N���@��!��
�Q{�1���D#�C��^�5�DwL�����}�Hu7��v�`oH!�x�i�t�a�a��A&�']��T��0�i�8Kb���%��7����Y}m6wGh�@�$��Ź��d�Fo�X({�5<������[���!�̻�`��l~\���|�l���}�c��,�!�����O�٧��������PK   *V�TD�98- Cz /   images/ac84e508-e9ae-4a97-a513-a57c89513e93.jpg�wxI�&*�s69�l�Zj�e�b����"Jj�Vj� Cr0�`2�&ۄ�!�&�!��M������v�>�����:]}��s���ޣǥ/���"�!)--�4$�"}��$\vI&#e�H�j�����
)�S��d�T1���<��H�S���׏o6US6���}ӫ��>�5��&�"�5'U����WJk�^+��w��Ui����7J��RzV�����T��������Z~ï�:�K"�7n��O/ʥ\ʥ\ʥ\���Lѻ�X ��U:�@[��mi��4*�F�Ac�!	^��t%l޶��E�o�����
@�,*3�R��,�F"�G���xb���{�g��~�w��[H������ӦW��	5�L���>~z��XW������Mo�~Fڟ�U�H�N#����-���>�ʮ�w���J�ǳ+�ms>���������]��^/�����n��o>T�@��=�_z�?���bLuߒ�ޒ
���%�a�K*���>Y����c�����v���F�U��^�/?��*�o����/�j�ҫ�K��/�ֿ���y�jy�ozFJ��+�i�zM9+-�r)�r)�r�?]�Hu��Rʆ����ʢ���&�ՑS�J���$R��vR�E���˯R�_�1���~�o�W�7�oL�N��b�z�Z�>[�ܖу�|m�Z���������+�8V�5�D���V|���w����G�}��/Nv+��_6Hr�
��6���I'�Z}�����bS������A������,�d�Yߑ����z���2�{�������˴�xd������f����hVH����G*T�Ko[�w�w�o�K_��x�jU�T�R�ZժU�W�V�V�ڵj֬լAú�Z5oӺU�-�v�ѹmF��-[vau�F�1�6�ٽ!�W:��HZ���kլմv�@����i��+�~��g?VLkG�P?�b��/�ImR^VN�&?!*V�\�j��5j�
R�+�b�
�*V�\)l�_�J�+7hG�Ti�2W�5~���Z{��=������57iڬy�N��t�d�L����BX����No0�����p��x$�'���1c��4~��왳rfϙ;/w��+W�^�v��m���w�ݷ���C��={������._������J�?x����W�ߔ�}���׸RYC�_�ߍ+�^�U�T�b��_�J��jP�R�v�*8���P���j��3�n�S�=}�n	��Ѹ㷎/���-��Z`���"�;��B�U1�֯X�ԗ�j on΅k3[�,�Ж]a�����������7�Vl��HR�{aن��/���x,���7�x̶9Ϧ�eO/Ѻ���������Z����`��ꇋ�����U�5UXitg����z��S�Q�i��C����۞��fa�U���U��Z߷^O�i�첋����ϖ"��t_~r���m{ܫu���sk7�Go�Fj�ߥ�,�{��f�{����u��9�=*~8�u����p�X�f٭_{~!%>G�$z�r/�g�o�b��֛*�.h+��jm������O�~;���~���^���=��U�-}ނ?��O�������8�뚤t�)�N��z��YP}������w�r��~����޿����xڿ�q�iaZ�+�b�qS[�睇>���p��֏b���!��.ҳ+wF����a��Ht�[mpw�4�P�{�3�=�Um�`�rב;����N�ǚX{�SF�+et��]���X�7�=[FԄ~{��z�j���b����ʭ�]��b͹����t����F������u�v�U��v#s���]�NL>�k����ֹ[���m�G*�Ҟ�j�~J��жM\}���J�:�Kmӣ�y��Vx�H�\�ҷ��ͺ�|!��W���4_W��lX���K�/�W����jBS�������N����������¾���h@��;��Y����W~��_���7�x�8��mX�[�m���ٲ��Z�V$ON+�j�?�ې������ז�6�.Sד���?������,>����gY��>رܝ�!�o�R�tn�mg6읝ݫ�l�էu=i|��YiU?�ߘ�l�y�}�2�{�����W]q�^Ǯ��)3�L%����`s7_-,���o�����J��A����Ng���K����q���o��T%^��Bz��{<�[ՙ�f�}�����Kʽ��E�m��Oh�]P꺝�d:@>����� ��m<�sOҊ����^ �J���	��矾��:"�K揜5�ٻ���k�N��E?Qk�ͨv�B�Hv�۱=�?z�����y�/\5�V^�>��JyдR����z����N���+�n�q~ syPs�	�+P����Y�)�c�wl��jx6-�~�3���g�|¿�v���=�n��V�k���kl�V�օ�M��(����i&�m܅�p�-�tl[v����?�������:�iΕ!C77~i`�p�JbI���+�W�+k�3
��^��,����`�;3�^RX=����i�ω��.7'���֫���Z������r��Y��]�X���_H�lk����kscY��N��8ݱ�D���B��s�C�:�����c+�����p~��#�w7�+]�r�X���ᖼq����(/�Z�]�:`��r>?�k���OO|4V\!������KO��A�cy�靉W��7n���3�&^�,�,Z��N+z�芵��p�v�G��+��K���;�w���_H?;׳����6x��-���=�#o��P�(�@��z��va�٤���.���������{�NWaN�*�{5�XZ�F��/��v =���ӵ�8_���pp�5�7ygo�V�SKX�v�^��v�������+�M��-�Y�{����0�;0H��b�w�ܧy�{��kU��4���כ����\���gg����y{�i���`B�-�rT&���h�vy@���^�.�X܆ӿY�Ô�G�שƮT���m�����8}�y�,���֬�3��]y�kό���͌��M��S���/$�E���+�q{�����V�z��ΞQ׊%���cֻ3�F��24�޸Yڑ_��{����lo.���1�j�)��N�\g��y=����9�'�(�M���T9g���^����ߣ�1�;4\��H�q��c޼v�V���|!�>Z��ޣw.�F� O�Ohث y[Ԫgn^�G��|��|��d�l�n�t��O%�Qu�0��w��ny;tW�]��CIÙ�-�Fw��g�}���
�������#ӗ,_~��N�ٗ%��l�\Z��p�����bM����"�)|�8��:\�Yt��j� ��}�Ǿ��}Z�j!r���������s�d�k�KG��7�s���/�S6�cX:��㓴QmFw�o�r�`��m$�^���<���J3�?g>�R��-x����.QJ'd�����ӧW]%>���z�����ִ^�~��y���I*�-�"�Z�.4����g=�|>��Wc̳[�����*;��:��nO�'�۾͟6�|���t�}�,-z��f�����x?��͛��X8�u���/)�2�����u�ҡcx�s��wO�\o���q����쏞��΅Y�^�-m����(3��6gt��˞!e�F��7�Lν��m�k�]�����yJ ku��f��E+w��i�p
=�G������PQ �{�Ěۤ��Q�xߝ����_�O�V����+�y�o�(���������Ӭn�\;:�ac�������j�1s��v�2kv#M���������;�6���Lǯ�]9Kk=�"k�ia�3E�v���w�,ިqj��{�k���㍦%e�yK�%���**�H]N|��Lؠ[��:������Q���X���7�{��v����]Z�?���{��q/����
�8�[oV���u��UXu���;������t��ͻs�}�׃��)��|w��b7]8a�˺�e\W����/�_���u}pk�GH�d��I��ys���v���y�ǋ\�B<�7|�ԏ�Pui���G��ڎ�.�y|����F��+����ٝ�Z�b���o=��4ۙ?t���3Zι�b�q̢M;H�.9ٵ���u���-�
��? t���H�s'�t�Q|���A��̵��3����(}���7ײwduɻ>��`Wm��s��WG�k�B�vZ��K��%W��ł��I鄩;�e؛%<��)*Tw��T�V�3��b��-f����g��)+4��<X���4Y����xh���6}��Ã�V���SN�qA�mq|��׌ܲ�a�4�7b��zW/R�>6|�Fwҿf���n5ܐ��B���+l�u6f�1�� �%cv�'u�>5����ld���[[��e>�:xMͩ��?|�yr���6e=7򓧡
�H�3�6���cYM;KxS�Ɣ�.�z�<��]��>[�sG��7pV\m17�T]�:�b�-�����;a���~��iy>9{]h�.˰�i%�ֵ"�<<&i~���' y�4�l�Sޔ��,���ђ}��QG�o��%^�����Ck�i�ݜ3kWviP'�W�,Ž�ܳ�Z�͏/]�ݡ��6}��עUf�:G�=k"�^9ּ�H�*h��½I��RH�t�n��~�)�����g�a颜gݧ�_3���޺����[�(v/�^L��,oN�qI��Nq���ڸ60����s�3�5Ba`Ծ���m�ux�Ȧ��4��y��S����uf�@wlv��B���k�c��3o�*81t���p�޾ۚ5����{��{�Vd���Sn�񣤔ڶJU����KH���r�M�ꯝ��2����&�P��:a��L�jW���f����V%����Zu���Y��g����Hb_׶O�^x�K���n�gm����k�8.n�o;w��qc^6Rw��5m���/W����dH�D�+�k,:9�vs����_�4]�����a]�9�_{�4���|ͧ�puq�D%5�i[cp�5� �7kNY������s�v��ʭx|5W�yol1�;���_X��>v���;\���O�eC<��C~ov{��K����|��YݗSv�/�/�V�����+��t�����ئ6n��oiW=��[����%�z�Ý�L�gb��m�kl���;��b��p^����ת]h�l6�x���m��w�����r�1��鋟&j��"雞��o�aαs�V�x�;z|ݶa�k>r�v-�`qV-	�<�*n%���Q�'�~����SWըVa��{^�ӅM?�����G__9�W�&�{V3;��{������o�f�ޏ�_��hCJ�r,�7�dcf߳���Qr�X�ٿ�Zwe�U�G��S?ܺ&�w콑�h���A�z�s��t�������؋:_H9�~��9w#�"o�����,xr�CɑV�d�%����#];�� ����d��E^��d�q{�CK�.��T[j�x�K�p���������N���G->;1�[cBnq�]��3W�i3��'�ߙ�p�c��ݑa��sO^�m���S�a�ߍ��;��ҟ>6�꨸�g�7�c}n�8�k���&��Թ�N�}drΘ&�9��}e�즗�}(r윂���m�D���f'ZN���x~�5i!�[ր�f9�0"k�Ӛ�}��ۿ��[ȸe��������.ޥ�-�����yɀ�>�۷P������BS/�Oϙ����2%�7];N�륤
��}�������R�����Y�6�BQ�Z�N��/c�z��]�J^�@B�y[I�[������&T����,�ze�@� ���7�{�>m�s��Ӣ���;+�LXA��� *����>pU��w�s�+	�O���:*6��u��}|\銩�e�v�}���Uhb_����cS��N nC+����;CFx����V��Ѷ��'�W����|�|��c�b[QA��#�)����e���K��UG;�������]����y��?�r�ww87��[�Y�Rd�hĐ�rp���$?4�t5g����NBj��Xޚ��-�rsL��Vx�e��h������lQ����K�������Z�,GO��������G�MT��_�w�����<ٲ�sl��j��oZ4ht��ѿ9ip��ؚ�?���tn����ҒG��S�)��r��ܤ��f�GGO��sЈ�}�(�f���m�>��څ��ؗ�n�ԟDX���l"[;�V�3�j�����璦~�T��UГnXF������N�xz>����^6p�~�m0�������3w���CG7o�x5�H�i��q���۾�ށVE�vU��)�����]{W����~�K�3��5�`q��٤:2o���vߧ��?'�|!;c��¸h��D�C^���'_ߺ8���6Eg|���}�?�h��|��Z������6��k����=��է�d��ݺ,V���ӿ��.N!=��������_�8�NX꾓�?�Y�d��jS�Yaߣ�	���=���a�Ŧ�iĜ��}̭�S��JS���&��#č��9M�W\�ƌ�5�J}���xe���ú��_�b��gZ.��b�u�|i����Be�״lHv�m�Z��E%�~�;w�ѓ�?��3�m�{^��z�xu��i�{ͭ�ы?��������,�:2��{�OF�Lʪ�S(p���J�}�jЪe	Xq�Ž~[DYG�Y��7���p��?X�r>��Ǘ���ʫ?`��Ȭ\v�ՙw��~y���������5��ߦ����?~��9ځϓ>o�V�����]����W�e���h���L�!s��9�������d]zҎX4���vIɵm����j���^H�ʶ�$N�p'��5 ��d)z����F�����m=�>��ο<��akŭR;��by=#�-�e����\æ�	�km<��r����n� p���B���)j���'mg|��͓��<8e��ꕞ�-��������nE�?�\ś��[j8=D��z*�!~fhu}xvs��5ޗ콫�0�^]���O�:�ѷ�m�w�؏'k�m�~F�*̳��ڔ�S�F���ͳJ38�'�7˲{5i\����k�Ͼ�H9qצ�'�%����ΪZ��n���~Zk�Ȋ��n��]�k:zp���f_��]P?�yh1�x��};۝�?u�:l���O��Yu��X:l�ƕ�,e���N>~|���C�����l_�w��i���M��Ч`���W�"�_Cw�ͫtџ;�3:xvQ�N�CC�>p��&%��캜#zD>��w����VQ�w>zbѨm+Z����׻�V`$e���H��D��A�Ot}Q���[�e:)m���o���G6�5m�"t����'���i��K���;mv���\��ɯ=���]9�n�k9�eH�{=�����[w�[�}'S��,,�|���|N񫼛Y8�Mݢ��*��M������X�r4qh�����}��;�]��B���8a��7+ݬX�N�����i}���}��)��K6�[������z�B{z��3��B�N�G�l�szMC��A�O�����D�{���4>�p��%��L���mG|���.��G�qF^?`S�C�,ʥ+���<�r_0ĝ(������t?X"5�B3�q4 �4�le�?������닢]�m��bn�>��������X?�O�
[�%�ª/�w+c�hQ�s���]捳�d�(ޝ߱rE�B�����j�����W~!%ft:ez�_͛�uLnа���'�[�Ϟ��cS�D�99���6@��+���I�7Qefsux5���
�G:���$>�}vp��3&.����ר��o�מ:�>[��!ZM����( [���ˋ����-K�oUu�c�S�����c��?�h��:cָ�u2l��Z��t����f~��І��[d�F>���2�?�8���r{��Ⱦr�r��C��/,)�1�V�;�\�{�yخ�lQ�y��U���ߏF�����=��r�|�b���L�)<0th�����;���>8)�J~��+�5jpb$~��U-���2����բ��@���0.��Q@t:�n�M��ir�S��{�m/���Z�!p��ԣ<~��Wm�m�VڇX_M�m��=�;������-MX���ǳ�&�^*�p�,n�k�)�<z�|j�~�ҝR��).�Q l(zz^��y���Q﮶4?�{V��>凉�l5��(k����pT���!�Snux���(p�v!��y���#2���}b�Ӊ[�4��Z2*�Ҵ��О�����pvN��B�7y��ij��z۟�z��m׳��{�e�`L}��"�}3ǫ�M3��\�����r;�m{=�Ɣm[��/z8 S6s?��tj�C���j
�$]��|���~G��%�ۣ�:T�z�����j/��{z�P8ᘟv���VU���mݙͧ���!��?j�(˙��-*�{�����Խ����
ۓ��_Hm�T���w�׮�s3�d��Z��;���z��ԇ�����<��ǟS���(��P�a h<��WYO���vZ����iϴ���+���?ɊG?�$�;�䒖�n�-�Z r��k�ɚm.(�p���ݲ���*�
g؂*}�S{�?9R��w�I9�,��|������$�V��[���R��MoZu��z��mu�I��o3~���#�[~�����5��S�&�\��9m��^��5����_��@���Q^��P�Y���a�<���*��T�\:�,�7)g��Njz�Z2��<�݇��^���Vὸz~D����`I�A��O�R�-0R|��6��;�\sa��Ntâ��6�u�r'D�-�6��v�Z]�(.[�*��ؙ-�o�����ȋ�?��يLc�v����&CG�uN�B��wa��T��V�yW[�`3�	��G�>�KYZ�{��鸲Ik�����\��i;p�ě��rY�g���rݪ9�Oج��� �tc�w ��.��`�hU�ة�����)P���x���f_�z�s{�*NOw�H�|�Y̓g��7��&?M��`���7nT�u��A->�dj����޺�̫D�]���QG�L'���g\|6��z���a.Z�~���F����U�T-ٜ>� ,�M��7��m���W�Z_f�{�{�����g��u��lWG����C�t+�w_k�Ay��kЮЉ�%��?�u|��:�=ؤքί�m��}rw�{���C',�O�\���{���n������`W�/g^c��ޢ���g�Ϟ�vƽ����+�+�r/�F�چ�'��<?�j�c��[n�r�em&W����5�����5�<�^O�>�^�U���<��u�ܪ����H��f��Dp����;��{��U��[�\���3	fQ(~��Xl=�%aRh=�R�DV���"�	�׏g%zg|3�J�_�)m��D<�38_O�5Ȕmy���-�#�Dw��J�g��]�z�0f�B���-��zg|���=�����Bc��*@��)��8Ꮨ��x�om��߆[î`���zl��������߭�������W�����qA"b�c6,�|����r!!��d@�ɢҙl>�1yL@H��ߕ�����;5�O��M/l3GaM ���_���^�����?\�^��䔇)��n^���RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR�'��&�f��ik�c�;�;���已���-��"pW�O!��m� ��V}������������+���7��ݩB��o?����o����K�_7f�߶o�������~]���[��m�Z���i���E~�M��5B��lc�	D�"�Pz��B��F2��a.�-Ґ7��	>[H��B��F	+;�8Y�T����\F���z�Oc�Q�^�{�	W�+8L�4F��HW驘��B�b;Y�M�cVvě4��	�Ńj��%E��
((�����N&�b�,�j�\�u4=*r$��9iLI���`X�<H'cZ����)��y<���t
�C��ð�a�+)P��ܐ�G@=n�|��-ѲD�Y��%XQ7K��Ǽ��	1�

A'Gȸ�C����P$��D��#�j�`�CZ����+`'�I��]�r�^?$���J��k-����P�W��a)\_��D�Ŵ��X�N��iì�AQ��ƹ�hB��l<��œ;�㐨Yt�L�cQ��8%��|����@1I�/(��Ȑ�m��bV��7q1=`)�˙	��b�J(H0Ĉ�p����wLQ8p(��'d��`�X���	��'�x�ڨ\!=f�� CǑXT��=�&���<r����Cnf�th#N��o�)MB2��:<�^�Q;b3�uv�2ƒ�Z�U
���Fx8 Ć-����F@V���x�+7r�r�SF �@�rƽQ�U��*��!���l��J�	�^&�Ài���g�'itn�'��!�A+	�"� 90�"�9�lp��[ ȘIU	��44��p�\��d$�r�e���)��vȬ�Pe���W�ԀާQH�Ar�,ǂ<��k�[ �h�#�<)R�b���i��ԋ�����q",Q�>�(ruj��	����>6��P 5��S�^���ǵ��w��4��a�Z��N��<�0bV�@���{���A�{z�.°D�
��qs�zq�꤄Y	�phh����h�CD-��d6&��d�5�:|.�@�d��,v�±�j *`�4��e�Q(�c��r;%�R���+@V����J����mb;N|y��s��Ӹf���)�jM
���_�Tv���D�^I�eu�j}.=���<�E�gQX�$���f����)ƨ�$�1����^V �dFMD��*����h�)�bW��
`6����+�X�$�N�?`�a&�mb���J�tI�BǥR�l��z��⇽QZ��Q�:@��ZEK��c1���[�DRn��0A��ҭ�ek��]�y���
<4��.g��7��N~���!.JW��q�]n&b��OE� �0RIjQy	mB�A���*���)���f�����2���%+3f�1�qyg;�q16���Hjx�!#�&q�,S�Z4 ����o7Sl��[���[�z<�%%�7 s�N��*W�a߬��1m�́y�3hd�ɺ�OC��� Kb�I,.[�5�]l�:�Ǭ4	��Ƚ� U'�����yr���T��(�2� ]��n�)�Bv�
y(:�U�#��+G�RC���:�'0XQ�֟�/Xh�8��1�1�l:����C L0�̈�
KBoǹBN�+ ,b�G�{5JwBI*��#q�I��*�[c2�KB[U���Aj��(��̓�J}�F5G��8#����-"7[q���"�iW��[��L|jHm�re�����Z�Z�	�U�vC\9��)1�����d<�!��Ef�K�T��. �P�u�%,�#���ju#:����0YF�B�U�a=D�I,q-���lB�Q�4���s�5l(d��T<��a&�� [ln����(t�Ea8�^zҠ��0�0#��.`�D:�N'��q+�j�[RC�@�7�CR��&��U�Bh&KL�&�Y�
C����.2��\�ʃ���(����Z�P/$��@4�ٓ���Q1�zfR�Ty�����>)��
�sʓt�[��ˑ(��%�� 7,����Fֻ�z�Q�\Vs��E��䆘����Z
6ْ
��LQD$r���D4n5�+-" ɶJܠ��" \  `�B��*�O$�*.��"I��H�gj���"&� �@�7��-�YpS�)f��,�z�9�
h�?š��S� XF��I�^�P�h�U�2T�`��̐T��L;����~VjT���@�b׊�$K(��^D�� W��b!�)�3q+�&e���%hd�:g��|�6��!����]J�Id
%�&3���y�J�b 4az�A��@ք"�r�Bc̭���Q���*����A�Q3��p�f�$����;� �c�j�?�E@9aa	r�T�%�p\̶YWB�p\@�Nm�%`qTńC��W�	Yh��B�Q�A����AM�ƨA����\I	#,��6W
3(5�d�4�֪SDa�A���D��J��L����u ���,y$���S��	M< �C(`v����Y8V�p�U<�1�%J�GG�IF�HfƜ`R)G�AJH�y�@ܤҨBZ6�~�,��R��fK50Y�s�I%, h��j�H8�uR�3ƖKQX!�@+��04�^�5$�HM7c~�A�]��Ô<�H,@�q�����E4�Ӈ�5,��X����[uVjjf�KD�W�ԃd9��������*4$�'y�U.�1�B�����R��͢�q�Bfa.��j�x1�q��&>ǧ�m!�9bV�02�"�PB��F\�J��d�0�r�9�P�|&�)*#		�<b�h�9��6"΄�h���Snz�ހ֜�i�>�&�Q=��Y[�+ӒR�FX�l�N��q�:��/P�to��І���)�Z��ēR	9�K�2_Rk�X��0��%G0�<.e fr�%�g{hr��S����l�s�e�T�&�#	
7$�q-��+����Ԡ�L~�(��J���CAE\"1_���MR2O�
����9��'�H�d��k�*�HX��E~�-�Rm�0����� ��G��N�ƅ��F��Ƹ]�s���w��J����Z�UP��f������;�*D"NP�@2��+��V*�QSO��i��H�=����f8�Q���ѐOY��<��T4'�d�9��J�ɄW�p��#"��I��pȞ��L����N;M�	C��B���<a��*i��@&�c&.I%W��.�CV���7˥R[�Ű����!8hv	1L+�l#F� �uz6;E�x� ǠgriF'���1���ƨ��-��C���m� }��0]9�t �V�I�4�J�h�3"QB��^eN���0�z��S2AXk�I����ϐ�l�0�G�L������TK�j��̴�-&�1��flZP�5H	�N,L�N�`�nD(�����d����&�G��ڴ������ �(Bq=���e�  -Э
��	l�%U\�5�V�F�4���*��
��L�C
�l!�/��,<�Ѹ� !���D��FxF�h�d����Z���,A�
5�<	���k�!=�G(�����U�"Q��L��bp1&�d� y����>��A,@06��2�2�\
��`��d�ht|���x0��ń,"E*������c��FĚ������e!���
��1qLtF�|D)�"#�~ 0�Ѡ��:�����섣�_ǅX1~@��S�K��@L�Z�MV�&��RK��l:S���F'=:V��'Ry>�`̑L��F�g��X�e�d�V�(�6�0-��B��1\j�p$|�q�mN���5�%�TW2� �3�-���n6�/�H����)@�M�A��J�}n�>����,���YBfk�)t����0'�17�E�bEwrur�ŭ��H<�j5a�ǝ���-���"�t��j�r'ZJ�Þ�0�tr�V�]����˱ ɤCM�a��/O�6=�G�8h4�Sy��'��\(�aJx(E�)I�D)6�L�+l��C��G�.]��`3���ð�5�P�JM�Hn�3؍B��nv$T>TcZ=.���X��ː{SD�	�Q_�f��SYM�|&� !R�|�Q���,y��BP�`��{�$���LbK�\|
��I*���L"(�rj�р55�)Y\��(P�1]$5#f?f�Cx܅���L�,��J�cHT�sڅ2�����I�9�d'|V��#EBS�.������
����vS �m��;���h(1�N�Q9r�3�t�
�&`^"!�D�\�K�TSL
�Y���62,�1S�{,"V)�����0�[�7Q����d�(G���;iH�	$�r��K�S"��M�S�K�D�X��	<n/䎲�N�����h�88t3��}��BL�RJ�
i�j����RO����,�*�Ѡ*5��0-� L�����È��V3z��f�c�eLPx��mS'�T}05��cX�Q[(�>;/$�@�����&���2�<5R��M�0�"V��	�*��E� _�F���AL���N
�1@a�a��TNLG�� �̠�L�[F�6����L�U�M���S�M NX�J�	uĸ�΃%D2<Lh=4�COXi+��(�c�KĐ�$��H�F�Pb�#L:�F�R���6�FC��l\.��hF![�"�̨�i��V�n�l=
Qj�C���-ۢ��27���N�¦�P"�	�.�Uz���}ى��!��)�p�R��L|�cV.���6+�к���M�Kz�x�M��Ƥ��h�K7��4�����L:�-J�r"�D@!3ðQ�b�	�	��:��DM2D73SY�ܑb��0C�kmj�����4�Io�'6�-,�GM�K�R#n$�Բq�K"&A2 J*!�>$�蔈ˬ�I�pBLn�DR��09t ����1�ˠ��l0�)#����B:��8�\��ة�AMe8�;,C< ��h
Cr�-�yi|��*�Iw:u��՜Te�%����a��̶0?�2 �de�j\e�1.����>�Iq��1��PŠҮ��:�Y������&\oԅc~>Sᷢr�>n�sR�6Ȏ��u�ꂩ����-�-�!\�g���M�J5�*��F6sX^�r�v�������]��v0� [�` �W����̘+��S0 �����%!�2G�rD˷	�j�qDa~<ŗ�0�.$�*�/�ƃL�Ds�8=���),WF3�f?�%D� ��) �oS�"Y�P����!�U#�b"@�P�|�o�%),��D�4��*�C1&=��S,�H�4(�NA	�#Ŝ,-Ů���� W��q�	�SSc��b,��a4P��P4��A=_gEd�2B�����v��!�M��v��g�2��%�y+�b�4?A\Q�'0��CZ2Y����W��Q�+NUzV�ȄS�����r�
V �a,�_�Q�j�3�|��t����NM �T�T�BF=��#�ٕ�������q��A&�\*a{:�A i&��oF�L��W�A��n	��B�b?��4a	�Ďm1�M���Ħ@��SzA7�#��c1+#~�E��I�ȉS�6M$��E�`%�TFj���1O܇�~���8��H|N�cz1K���)v�r�S�4~��I	RM��e��4ɘ���P���0H��>y1Hc���,�R�H��dVء	�X<	� �թ�,@T�$�0�#�h�-�q+U�B���[%�Z�h��L�����HjEÁ8Yh�@qa��b}*��?%�D���;��R�p�#r�_%�Gck�,)PĒ��	3�����*l� /(��2!᪕�`HOx� le���H��7�dl�>�W�ZT���ܦ��L�=č���z?U"��L:X����V���'�:-9�'S$����E�]
� #�*r:]������iI2����DJhYS�a��Ga��x*�;�<a"�dX8��? �
��t>� $Xȭ��$,E2�"��a�D���X�4�ۨ�CI��`�ͼ�\�MX�):OV�M��U봘�Ǖ+@�����"�C!�A6��Έ,1He�bZ�4�ē<�D.���_��-��F��4I�%�� 
,�uQm@g�d�8��@(!�H#���N�&ss}BY�%iat�&�Gav��j<��jq�̑�$
6�a
؈U���S�𳒩�ɅኘY��ꢨ���,�5Id6���$T��PY�VJMP�k�ʢd�����*���I=�V[��vf)�q�q�(�c^�8�!q���B"����� ��4�E�^m����,�$��(� �q'q����T'��{��)z�)���`��_%�Iƹ�
��@���S����b^���\}�4rΓ�K��	W�ZR����
��
�'�ϻ2�X��K����)�R���~E�M�g���mL-<���N$Q��j
�
Z`��[l�a�ze(}9�L1*���c���
1�D�H�j���]j�J�p�q�@v���,�E�3}v��+��"4e�:�o\�q�^G��Qi�n�L��/�Q� b}ֻmw�4=`�W`S��?{�3�$r K��,;��@��3��`ʫ����u�H�-+��dRqcoN8n��@�m����R�2���������b6�p�s�A{H�m�7dݴ�;WiL&�ǖ�걍R0Tm:�iK���?���7f�c���S�y�*���35��:yd�{��Q�=�M)�-~�ƴCk��y!�Z�T��/5Q0Vb�2E`����^D\��H(/|� �ry>�\tN3H:3f�P21v�i�0�mW�+m����B��q�YM�����L&��8�����OL�!��N�Ĵ������+��E����]+��B���2�2��vY�	:����	r�n�9i�1N	��Q�!�ЇrF�8n��u��[�Mx�ݺU[��x��ۉ�ϛ�����fʜ��m���
���ag��|���hbS%4����{0�d}�U�Ǥo���E�x7�	P {�f�
M�٦�Q#P'�@h����0`x�~�9���]ю�����%>������5�Z��D��+ؿ4��gl��:�*'G�^
��\+�3v0�c`OK��b���s���Z��Yg�o$9����Pb�f��6i����]����F��< ���Rn�(�B�7J���R�\�%���F{kc�t��X��7��&7XvG���pn����`5�:"��W8:�P��wW�QM&e�-�C��ћ�ē��X9!��Bپ�>Ѯ4��z��Lr�`��W`Ο�h�|δ;��E���n"��gM.1Q��T#��I��T�.�#�<`D�2���Ld�*�h���ha?G����X��>+��g���j��&\�8�� ɵ���o��N `�X��oFv�S�+޵�0Cd��O�?��zq�M�;:'�)$�^j?�{�^��@��,�]���M�`1_�������@�(�p>|Z��R�!�&`<D �FR���Ѿ1聡��֤��\��9���5kl��g?�n�P�l(�ק�[�=��%��!��4]Xi-��n]7�j7��3���	��0���M�(�
 ~�����lf�m��[�����3��E%��t��]�;E����V���Fgq1�+�E�S�?�Y6�~��|MW_;&�;�I�һ^��u��.A���9J�M��3پ��4r���:>'ƙ���rʟ�}�0�����x���W�@ݿĊ�ʾ,�zgA���czپ1�oz�"V�qGh�Et�jO%���0Zi	��M:�@.�y�^���M�
{�O��yuVT������F����ȵ/ʫfC�YI=�~1��a?:��*!j��8��,ϧ�9)�?��/��M$`t�X�#��W�IՑE]V���]�DX��śbҏU.u�+��� 7�yOC����oI�0j��Nna��]uC˺�	�;?Ɓb?!r�4��1M�~�~��U�ѹh�(x_U�a����gn����Wu��8��kzS�����%�r�p�o��M=�L>,1!�.�� ��<1ո�#�YiWs�!F	��T�@o|�e8�MY�#~v��3ٿe���Ҥ��`dN�^ �0�ތ��xq��a,:�-�Xh���f�	����|{� ���Fx�G�zZ.BN:sM � ��t�Z��� ��_5N�߇�}�E��^�
`)�?���KB��j!\1���f��n#������oD��ʱ;��V͋�Is�Xvz�p�J�c
r;�c��{R�����y��R|	�,z�-���	��tf���:�U��w:��3~��^�]4 e-����W3Je�$@}S|�c����H��f��:|B����w�����R���C�9�A��28����8/!��Sf���X1h��݉��d��D�s4gysŲ�y��:z{n^Cj�=m~E��'���J�z��0��Sua+wRA�
��ah>T9��P+�,��/Cw���i)W0�7�X��m��(�Y�s֤���R͝V��ld�� PJ6�'�
@&�[6�#ݝ���P��,wmB^�&}�F�2x��C" �� ���&?)W����u�_J=�蔆�������'���x�O#��7��L,�!'�9�������vA���sF �	�:XL=�y+�9�V}�58T��^�W�֥��K&�9B�ơpo�e^Z=���㌓;@��x��^���8��-����ZeD��<���*؏/��e �H�6�5�ra��c�e���[��cɕ�s�es�Ͽ�Bo�}b����`�3�9�������zkp�P �C[�\��9�O�=��)�/?�6�e���(��`:�c=���s��9ǽ�9FI�7(�s^R�x3�\���0m'ݻ�v1Y��哹�j�z��hg���%f�U[�oGN��)Ҷ�ܖ`D�C�G�ᇑ�g�����<#F<�WZҺ3]��&�?.p����5 �����w�8k���i3�	?�<sB�~�f,̤{����Ͼ���M����`ca��C"3Ҍ�>��{c修!�̅��j�B�m��4�l�_n�ϱ��ۚ�W�v�d(�A���V�'h�?V��R��n��O��&3��Q��\��sұ�0��#arέ�Ȑ@��%v�0���zj�K�P�޷|m�Mxj�/g�pDO5���6m�4By|!Tv���-�Q��[PO�{������k2.�݀�u%+b�� ~�\7IՌ]
<X���9n���T�E�3�
�]8keJ�ͦ���9�p"�!��$��LTh�Nŉ;J9mc�?�ո��׊6-�΢J�v�?ɗGZ/�_ńZ��ѹu#n z�h����C��)y=����g����� ��ٷ��ﴭ)ƏE�@��e\��.W�{0��N>kA����KT[C>�Y^�P�!�����o&�C/��@j3ѕ�s��},5M�g��Ֆ�\u���.��� �ƣ\ ��^�d֗�%,ӣv�׼֤0�dPP/���k$�0p�b0r�p�����ؗJ)���=S���W(uPs�>ѥ<����s�踂1�T��;���� �����J�[�9�v�Μs۩�!�t�z,A�l��┈�YcRV�,N��3=[��ŦX�H��IL2'(�������.��,��Ox��|K ����hN�V�@��e��')0t�vfw�v#����t�t���$[�����t&�1����Zf ؈�;���Nq�_E�v��T;q��	�����ޖ
�-�]�Q<�끪�#���Pt�U���bmnl+M��tT��Ք��tL��l�	v��b<�L� $C��I5��`�1�Ļ�����-���Д���l��-E��������v���;y�D�C¯T��y�� ��7!�����WJ�6a�[��S��������9;MA�>�܇G���-$�;�t�\n�k�O��'�l5�L��?��l�ٸ��l�k�G�S�LoAnL.j爞��1x8�h?+��V�(wn5��,��ߤ��}��c+��>I�b��N�U9�d�d����Fb��F��]E�e�<�	�����[�)`ꨒ�Z���C�C��@wn
"U��u0N��M��q-Z�ܲl�֗�o�`�&z�s�赻����f�����h�����
��>�50
���YE7��1|mR�d
�v�qE�b\� ��IG��O`6�:;a��1�����}~$ɏT�K@��/�V��@��&N��!�`���DWK�X+BRa	�0��1���s_\w�*
ŴeW�+3چ�g�7w_m��M�\,�,2�t��m(c<��2���wX�2]yسkG���t���]8��z� ����!�I�����*o��в�7�)��#Q��)�y���0�W�6$�����ݷ�>m"��6.ݩdsYu��Sٿ�$���{'��\nv��ʠ'ry�P�~���	�������3񨔣��A�w������E�
�7�Z-� /.��ظ�!��!&T���sMu���1fvaB�OJ��r�Z����uN�S�㍫��i�bf��(#i �+�cQUn�a��NW�z%о���0XN������W�@X>�����Le���N�ΐ�-XNqZ���?R���I��̑1#��ӱ�s�j���G�sn�������ݸ���cA�)��ڝ7���l�o�����~Κ�!o���)\��������� �߂�ޘ��sq�O��	P�M�k5!��F����.�LN��}��wm~M�+y|���4=�=@�1����@��k�kF��LQ��Z��*�L{�:��a���!�����u�d��b��������۪��6�l��\OjoC���X�&���>�tV {mD�G����~��!<�����p|[�����>O���2�A�)	�9�;��2���:��?*���W�����lq�����5�Ϟ���<����N�`�0:wd~��b��}���#G����~�c�ϏM㖔c�p�hx֒������ćI�5#�f�`���ۿ"���$Z~���vr���D��s��V!	B���&3`NhՀ�zJ��B����.�&Fo���H�|A�<5�u���D��0����P7ˊek|�b�_A�h��֊q�/
�FɌ���f��!��M>^R�9^����у�0��ض��x�@ô����l�_-�>����DaU�g�R^�������� ~����K/"ס-�F���*�eoW��_=K���e��KY����	���~�,�Ic ��<e�e>F���Z�vöa�������ΰ�sM�>��	)�"���<ok] a��.^hd�j�"���T!�!��Ι[x]�ؼ]�ؠ�F��h;��]�,���Y�O��F�� d�&����m��N�̾�$jj٢'��D-�@2
9���>�&/s��,ʕ�d+L� %W�4�q�b��R4�-k��80����c#�Y~��3�ژ�y�=�Ux
|���R	u�E�$x�fn��џ9���B1�ج<�gJ�H��u�����owpM��B�{����K��鎫���D�%�o�r�Ɖ�dj�[�C	kM�]�����c��>�s����;��qї���i
W��R�A�L���RK��f���$���kXe�v�b3H���T���)ŜGP�o5 ����vU�����c%b����j�S��s��kTa}�N��ʰ������c^��]�4�h�[w��[=�vZ�LӬ)��~鴥�����[����ٷ�`e��Kzy�SP�>��,!/��-�'<��ʢ'N�]��as��m�4H��*�1Vd f�����>�������H�2�<e�_��s��؂��رAK߷:���5����=mJ'�CDvR�Ȑy�WT��qm��??�b|��/��ƒ"7�h]�����)y(��t��8�ag&H@�R��6[�L�dsaZ	��7і�nL�(� PC4B���P#w����h鼖�G���P���1��vV.ހ�yu�0KP�AQlJ�155���E�F�N�#���_ĥ/v[hI�ǚ���?SdG1�\p&1=aX�!z����_ŋ����l�Dx}���p�=��q��j+��5�l�}�ͭ���
oj�Hpk#%K�ع~��HV�����<�g�|��ĳ�/�����N�
�.]��c�7#�z@*�n*�k�PW����e|�1~��!6��3Sl0��/y����jdz�9}R�@�F�˺\�Q�++�3b���0�!NsGǠ0;~K_t`p2�	!�g#KE]��
g��?U޽_�O�{�h���$�w�h5���Kvk�9�@]�vpm���T��X�u{������@�����q��>7p�0<A��sr�6�rN���6��Ub����G��}��oc�+#b:1����~�̐�>1�-7���L]���;k���n �=�"#�re7 0 ��7C}v"	'	���yP�_8d�sOy����o%��VW]	(�򗗝t�B���4M�b����0X��M�	�<����7�|E��$��H3��W}��Pk4�&�N�jzR%:V>��r������>n?�F�r�)F*���J>a�Ȑ��xz�]�v�}E�'���_�^V�&m�����o�;{�岅YZ�N�FvTSz�QGX���K���Ԍ%������?�Y�2�K?"�����KS�W{���;��O���4���<m�,6�9۵/N=��.�kt��2,�S<fT+�;����墳��n�䝩�*��I	�fX�~2�#h�Њ� �Rk*���I!��>S��)��*p ��C,NQ��t��E �Q���.[��<w����t���+�`|�fm�&�}��� ̰��`	�vy��s�ꕲVN��kf�<�
�D8o�h�H0Ra�gK�~��!�uh����&V�U0EN#-���c]Τ��+�,d�g��OgT\���6��E���Y�[G�#�s<�ø h;C��������9���$ ����`�7�O�����n�:}��Q����i�A�S��.Q��5%�r��t�i/���V>(�"}M���_4eJ���XJ���ЗK�ݝu~��u��yjdØ���i�>���-���7���#e�L�b��s	�JPL)�N�f�N:�I�P���p`js�V����ޒ��D�˔_�?/�]{��;ߊD����%�����~ ����]G;F� ɗn�՝Y8BЃ�1G�I��+��Vg,�%R_į���ǻ:@���9E�$T�`�?O��^V���8��ۿ��Ka2��I�&k5-��"�W13U"\Z����44�0����{c�O�,!߱�n2��A_�O���� � ����㫎K�n#˻�vX��m;����;.��З"&M���1��:W��8^4�8��0mLw�e�69�ۮ��
���kRv���/�F��e��9E��$����%�qWvƻ����/����0��Jb��&��F��-��~�����ae���0#�����M��z�usө���'n����� �}�´h��ލ��we�_�'Ɵ�BM)�����*�C?0#��/�K޺1|@�V1Y��h)�JF?�3Y�Y!��g��Go�nԖC��^@%����@�3f�����R�O�|s��d(A;\��,XPP���}a3�RU|k!�2���p�p�c,�m4�~"�!1��[z�k����1W��C��p�x2��^3%�ě[8�ssnK�4���x8��E>�����j�&�����O)�����SE�mY`�'�0�s+F��-@��/�9�B�f��> �%K�=|^ '�G��nM�&�+�U�����m�@�o���aq�iK[�nNj	�,��$`n7]��;b�kc�B��Z��'�}�ZA�b9Y�׸΄xs� [X�-��ey��a��5�;�׶�����T���Ẻ>����؜\#�ݩ�r�G#���[vM�S\�����UPJ�C|�S{�ߙN�DP�aى�r�HH-��5��}��>�����:
d� �$��%X����հ�a�b��q���!Zh �6I�g��ba��B��JB�XBC��P�f�n'>	yL��������&� ��@�?r��=x�a.����,wH?�1I��|'�qE��b!��Ȝ��O���+��o��cXK�ж�d����ը��R�4�P�8L�V�pz�P�R�+%^��Wb���r�q�J��NZ��Uk�4�'�s��`��\�b��i@�����k�O�~�_� ��q���?��P3x���u��!MS]T�-$(��(�A�=ߑ��b#&�PV*�΢���yź~�%��c���-1��q!��!�N!���\�ќ��F�w������w&�`�/�%I�������Z܁��:�DQD���n�&�������ι3��u��3�w�鋁�hZ�g�4��Y�Y�5n��-g�!���b�d8����*�V�X��D.g�,��a��(@�:L�"���Q,Ԧs��斎�@�'�;��5w�ۇ��p���0TG�f/������������Y���z�4I[π��*��.Ud+���Wq���B
ӱ��޷[�}qM8�l��.�)��Lx�=o�,�J�2V�%I>�&���(���"+Ӥ�^�3[n�����%0��3��Z/Ǭ�����#DK�؟/�i��J�+����*�˞K�|�"B���O�$H��b���g�)	j��]�"�Y}�t&*���[�\g����Ņs�
�#���#�6�I�ќ�|�/�S�m��]e�c8%c�)N`�I���_h����o�m���Ly
�9���{�S[~| x���<:aHr Ts!�s�(Y���I�"�fC8��\NR8�]:{�������1KF�Ƃ�q`z|;e����|8�g���y�n�(
Q�m�/:�N��`c��D3�q�ow͸���^�/,-rz�rK+��R%�|�ʟ˃�:Ŀ����t�]a�St�k+ejN��v=?��G,�9Q�e@[�0�)7ΑBB=틗�!4�ʧ�w
������I��S�h���#0�����C.���zii}�Tx�]�qؗ��Q�Q���3����ݫX��J=,�u�	%�4כ�I�Dw;��� �X����e|��aVK{WȢ��"�01ކ���v>sd�.��`1-rt���Q�}K�5����Tg[�8��7���/���joaiW�QȖʗA�j��InY��ђo���=�Rn����(��C�z��^�Z��(�D�V��T̴8���8Jj�}�:#~�|A�f�	/ƚ���iA�.���쪚x'^T����X��<{�ߞ,�Z@o�Ӫ�9��� ~!��+���D(*+
�s�@NȀ��'?d�"�2t���߷��~➈s[h%�[�0W�����H���8�r&�[������"+Xr���:���������-��i/���D�� k| �ԢTf�t�d��u<ma+�����>�D���"�^�yKQ�	����R���`
��\:���H6Ĳ�?���w�9gV(��v�fٞ���=s~&�	���:�M�Q��ݭ�s�w/K�G����V;m���Qy��]���"���t���Ț �M�(JS�z�z	L�̧(��wWd�|"p�ע]9L��m�
Ž�6Q���;�K��]�o9���S�l��?I�;3���d~�O��A�":[uC��ot�0+�PQ���K�3W���>�0r��ו�I#GlO��}�r���f���}�< ڧ�߷�Gæ�=�(�I��?gD9�Cd8Q.L� GH���Z��wZ^/*b��iՆ\�䂘4�@�LMI�jyv)�_��O�g���y�� ���Q��� ��n&rmK�zU2��.v��ě��Ze��Z��~���L��'�\������\�]�l)��8��_��2 ����k.3R������q1V�ga�" �z��������TlY=��Ȃ���Zi�g$�������y5�϶�#ǋ��  �xR!FCe��#%�&�t�@���w���e��ǆ�gI��5�*��1���:�
D����9%{>��_��MD�ZP��=�d�$��Z@n��֤�bT%#d�9�v�Ҿ�w���gٻ�{�y�k�$AP!��z�Ű٢�c�LcZ�?�^��Ew�]- �_~�6�8�gZ1+1��2rѶ&;�� ��U=l�ܑ?�Ϧ��G�x|7|����@x_MW����x��S҅��yo|+�]�p�c�0pq�R8�DIkJ�zPp��9��J1��.�L��i�ۿ��S�Td������q�Lz�j�h痈K�Չ�5 Z�a�fjA.��ء0�HZӗ�_��2o���`n�M���
.Um�d�/�;i��Ɗ�TD+a����E�I�!0%�7)=+�.-�O�"�-�C_�]�?�qB�f]��
��.6�����#�^LP�9�_g��_�o�uG
{[��*#��1�;!ԝ*w����h����'$�%�v�i_$�0晈b���Ό�|��REQ3N�z��b�7�@fޘ��γ�d��?�9�A�=p���)E��Q�X��<�|�`B��%�ԹiW����SR���|Ky�t>�a�$;�;��)���F�H�0����-�e<���\W[6�,\�S�|Ѽ����d�42.��X���|����Z��6��`�Y<�K�G�ySmK��Yzϱ���s$>�.�*����:<f���!��,���"�Q�5ִ���^����j�3��1P�����M�����i����<aG��Z&�#^��>��V�&�Jx�D3�߼
h*��}��v\�)F'�����+e�f�)�m%Y�K/��z��B�E��N�nͩ|�r�b��F \XX��	���m˞�(0��ׯ�)�d���Ө���J[}j"hb*w��Vsǰ� �&���l9�������#J� �%���V<�c��}f6����m�e~Jl��?��W>u1�,�����Á���[�ܭ�[^�
3#��h��%�׵����$�ά���g�:�i}!�����yG0�-�R��9&#}\��R>�z�Z�t\�h�.p2\��&�r!�
5��*Y�|�G�Nf��3@��91�4�O��~
�,��;�u����r߂a�gNf�l"����O��C�d�����P5�4����>���T�f�w��Z�AE���A^����l��_N�x�A��	����v ��U�u�rw`���2��Ě���!6��dā�E���l�y�G4�'g�]�����P+,6���
[�M��i�+��Tom����ݡp��h���[��>[����}���|��-�EK�鴍���.׉���,lj������Ϸ��"������+�^���gꉁ/�-�F[A�_�ԗ8J�W��1b�PD,��W�D�j��	rt]7!r���E�8������5���GvF����B�j.5�S�Q��u裌叔q�b:h���H.�︃n�����9���_�߯�2\�ւ?߲s*o�W$<�RbB
gb��i��"����O�XN�ԾV�O\<�����@�R�a�Rg��g����*�m�Ӷ�xo��.g���d*p��bʾ{���N�g�©���R�wwǹ����ò�������b��	k#�%���?�<��gK�XL���9o���q-�E >2����L�}�$qSW��L���ږ_�]����*��]cv�$���I%�P =��פ|�D��6�`���?}.�N{��z�ǟX�t��'�/L?��_.U����1�jT������V޾�S��y�
Vu�󾣙���h���~�]D�μօl�S�Gf�a$ L��]ℭ+�=)��5EP%ً�v0"]��2)������b��q��/�EA��vٹ��e�n����U�fe��u�#��:�2��;���q[��  kX�$�ҥȷ���_�D�>����͊;���n��h5������큿U��'_B"xA�<�!���]�17�LQ��#Q�'�̤\����x�\u����[�op";��ڪ�mr�Y�����b���$3A�K�C�\��3�}��?�`���ώ�#�� 6��ï8LY1��Ib�[�HG^�Ҩrd&������8;(��v�/�2�~��9ߺ���¥m?e�߃����t�q��戝/�bH��J�9W!�/~�TU'�Jx�I���U��J��e��2g��ew�Z*&�����PȰ��k�]J���%~�$�)}_���1�ԅ�	o�ŸY�� yK6Eܘ���W�Ұ���k�U���X1۾��i���D���f���
������o֦UR�-�=�k;�#>�=�NY7���x����YY~�>Ӯ�Jlp�H18��v��_�JɌ/0Jb���� ��*�'"Hw�v��%J���\+�ɳ��a����1�P|m��X������!&+����`����m{x�cr������ j��g��71M�H���w��DkO�k>׮����H��+<�4�n��@ϭ'X�<
iY	��ݟ�� �Ye���$�����F�?������ v?��RB3�������G�@G%�{V�@)q}E�	Ƌ�;ʎx4���-�XKG�e|wL�����*��.iM0̨�.�?���Z�Y&J?p잭��r)Ia|�B�	��L�p�Bҹ@���J�Q���}K~L���Zh3������+_[��䞯?��0�ڜ��-㢁��}q�F�8�5��Vk,I�Q���C���_U����1��q�
��z���-�b9��C|�
��:�Զ����,\�(� �q��d��;��鿀N��z�C���5����)H�]bt0��F�������kM�T��&H��G=�Ԕ8�q�C�y�r���O�y�>��� C���(X�? ��^���G&F�Z=��N�n�$�o�~"�<��ٓj�ؾ8C�k�f���F�k��;������*˂N�R�kf>����3%N��@,J��@�-� K=�;	8-�*v������/�_L���f�{LQxqR�s���:���B������X��I|yW2��hB6�(�|l5�C���W.����8G�K�rRO�ݑƯ����`m7����e��Y���t�V�q��ɟs�e��i���nM#&#��0#��&�53C���A��<������e�'E�G(��G����E9��vr _X��`�h��Z�{`觐!F^�L��n(8�x��C
9�����Rn-Nz@Z ~�������t3?�&�;�Eyz48*���EQH���ݰ[�Ϝ"Dw}�p�Z9o���^��#t��_�.����`�?� 4�r?�d����}��������"���#���v�С�a��ϙ�t2ȳ�t�<����<WP�!��j���s8#0+�����/k�Kp�.2uA��<o �P O���m.����f���Y���k
����쿧�1�82Sp@�CS�~׶[JПR���sw��� (�\8���:�mQ3�X��PM��\�l�������rxq<'�xO)��� `���I&�Fʏ$r��8�"D�	1z��a�yN�����^�]u���TĂ���#<`:t��*�/T��ŕ7���DT�X�������
M��|�2�Zƨ���"��4@���G_��d�&64�'�t���9�op��-+�?�~���2�= jj��i�H��P~E�U=ɫKAR��]���YW?8$��@�_�K����v�w�af�������Z�E�>&l��E�������بio�ކ$!\�Q��es	���t�^A�_R?~5�w��pFv�_������(LBkT�"#U<8U
����B�$�U�Bƺ��0[|vȓ�A��Ib�b���̘u��ž��O��#�I�~�_�z���تDh�뉔�$&�a (�6A� @����! ��� Ľ��[��yҹۆ��0�W��7�3lQv�$���+}Q�,�~T��5�(��;)���}����nCD�&bwūwg#} �$����	&�������^�^fKwl�٭�̟N>j'I#�+'�P\`�/.��=��7ӐE�`Z�)�F�ݗ
}ڌ�~�:�D��m��5d�e,�������C�/�vå����p�<>Ѽ�O�2*IЖ:���U����2�����F��9s�Z��f�,�N�$:��|������yйO�g��+�4�5uEZ��&�(�����C]���)�*�2�_�0�s]�!�A�i}���2��߹a��8ʕ�՛���4V�J�Qq�Z~!���0yz|=\��zU`8gH�uW9��ϲ�-Ah%� MdmH���Mt�_��Jr�V�Y�Rƃ���ݯ٠ꚉ5��ŉѭ�YS�Y��j؆�T������	dl��|'�zoѽ\�^�6��d�f���"�ҽ�tk�{�����/�{o0߂ �I�iA��l��Ɖ�@�v��N�C��rΪ~녴�Ax��נȵ�v�a�-����M�^���_��/x�%~#�6�0�8>*�W�e�Z�����4p�4�u8�O���;A�D���9!Z���m4<t�/JU��ڸoR�Є�f��z­?��kVe��v�V�ǵv�O�����$�]Ā�=��ac<7��{YB(H�q�d�G�N#i��3����za'�([P%�^V2ZT@n�3Эޅ�� %�R�e�t��y����Y��F��?U�d.]����:���.+\�䘞�~�� (V�	ḕ�Z�R���K�/L�9�֮m%Ň�u�8�R�Ҫc�8W��������]yc���<�Ab�W!����)��_5o��B�(xZ�9�!���P�N?�)���@�,���h`GJ]`i�)&�o��b��m�3�X�>JC����wqV��>+6,�t��k���x�sgH���� 7�0b�c��^1%@���_�<��P$$���w�ʍ��v'd��`̒��UUrΙ����!�Y�R;:��W��}�����U��%uH���},,d.��A,5w ꒩P �.Y*6DAf���{Gm�4(D�R���/��z�y�%p��'�&���n�@�ĉ��хM��������:��nsz��ت�6'p�[=}�լ��c�N��g��wae!��ؑ�P7��viB~N�|��Fu���9e�N� ~R��Zoݿ�{��O�I���bΈ��uEE�n�!�m���xW�鄮�{�{��#Źw�Ö]l��i��4.�O�"u�`�b�ŎQa�ʀ�Xf�C}`�4�a$-�;�dE�ئ ���k)L�����ϒ2H�⦕`�'�`���#A��at]F��aUsr �}�m�㏵�����6%���ANק՝t����F��������㵔�Ú鑐'8��n�<����?n�9;��AI�
�YrV��{�������n}���pN:�3��Ҙ���޵����|9l��?jһ��Q�q���o�|�q2�<�OviO���� �/z$V�{B�9Lq�pA�g ��b� ��R����;��(��QGJ}�	���(�4��nn"(b�5��x�ܶ�
�=0�>T��N>�!�w��5��u��G���\�ty�2	��r����q:��f%�
�K���gJE�
z�/Y���������+8�r���1N����"�2���U�֙�,�Myà���&kSv�t�R�xMzW�6�H �B+�{l,��|p7� emC'�>d��՛l4�$�a�N̟Uf�Gu�x<�]?ki1�ݦ�T[j:D[�2O�!����e�&b��m� i�͕i=ֺO�?�nx;�����bG�̾�^$qc��`�0����(̶Ӈ�V��B�+�V�/�K}���a$���t}�asIr{�����֑�cE�U� eHS|t��]ShiBB{��!����Zz�9��B��)�k��Y3� �&�׌�J������K*�`�������d�>
��,�j�O��R��h?������#����O�~� -_@֠�v���g�a[��|�Xy�ۅ������L�s�b�O�q*H�mֱ�U�"BW	�����[��kK٧��^��~�<� �E6��Ζ�]F �o�tΦ�{y�rɚ�ТP��*/�;Ƨ�D�'<\��	��,���87�ø=�O���:���q�D2�6_2�C�#�&ʢ0��bv��,q�D-�Z�7��X������`v?��	�N~~��:"�N�};�$��=�Јa�w%� ��/e{��?~���2}��@U��2�1�\�!���{'�`�w �b�[�W�5��g%�{{(������h+|�AH��،.�/&`��Xe{��2�D��V��8%FFerFܩb�@�Q�����\>����Ïo��¦���
�����a��f��U�ˁ��P.{�r�T��B3�1k�_ۄ�6��>�K	��
AF����mP|�Ɩ�1��XU�ku/�SL�A��`.���ӎ��u��X�����^��I�4\Vk����>ť��G��z��\P�y92�`Y���p�چ�6NkED�����|�y;b@ϒ��E��g�+�9�k5��+��"�	����J<�edݯ�����l��6b�YH�w҂#���������/��S�\ƴ�U<R�4#q�$D���n�X�68�Q�����i���ۙXη����Ɨw콉3����)ɆnF�Ճ�AYֻ��?�+��2e���v浾Q�������d��^�{t����Mr���<�Sd#s/fy����m�Fͫ�K�K���+�&�2��D^н5ݛ�|�8"3�]��1���6�6��'\����=��W���ij���s���Z6\��E6��u��I��6p���b�6��	z懮B�u\`���@�Ut�sW��_�^�qͣ���E�T:'�GD�Ym�R�'㯥ׁ@�l���:�>�чI6��ݎ�JKT�����:�i���4}�y��>O�6�_��&�M����"����&y���±����&gmZ��~�wg)NO�_M�efw��
�=̊��薒B�y��]1�zM��7e>:��Է�A��$V$�ĜF���2Q9h刁��:m�i����//��$(�zM���Kh��My��K�yu,m��ӱg/ �N*��Q�My���v�̔�S$0��L�s�f��k}�Ͳ#���y&����J����MԞ��q�#��$i�·��;�谘2��ޛoE�%g�������A>|�������b`3&���i��E-Qh45r�����>bjʚ��j����t_���B�����h#���XvK�5����$����x�pa��!,:�$�;� ePh��͔I�nL.��Le%��*:������^���%7�@�"g�Wwa��ޘ^���iH� :��\���kI>{�����gFz:g�",^@�`@�9 2:!�-+]��Z����_a��o�/�c(���7��#[�y�3�#2�@�|�x�+�m��~S�R@_�m,\"���l;]���w���v��Y��������8?�n��hvy1�Hޖs�%R�[1`�?����Ҕ0|���Ѻ�N���R����n�r��� Ic�#��v���qPo���5EbK����`����taPM��R}\E�B�솖�%Ә�עf>x1�[�Z�d�=�c��t������k��v#��Jp�c��5��y.3�
ع>��%��X!\�党z�;�`H���8ά�cE�t!�^���I�x1w�ïtU]��1�-�ˣ�4hn8��˔�����Ĭ8ѣ�p��f��@�\��img|�z�#Ί}�%=mŪs�p�|�6�RK|�J�D��o*��b�'@���}�c���K�";�9�oi��%��hBكγ�<���Gլ�6:�z��k��]\��.L� ���d��3�Y	��7���0~�v>�x����h*�'�l�;���c�b����'?�K�u��mRx�Vg��O�UaĤ�W�$qUfI��Q[�?˭H���l�N����y	�Y�!$n�P��r�j�a�bM��?�A�V�O^a�~ljn�M4�#�A��P�qD\�8or:�v�0�YgWja�2��E(��(W�c��E���
�_����_|������v܊k������!�*�hB��Һ)u;qz���9�t
�9�ly�J6����Ƞ�<��)CI�aR�7���i͹�t��?�v;-7���-�g�K��h�>��@������Y�O]�^6��w7��H\7=�[�J��/Wu�iK?b$|ܳCJ�/[(�����!��2�RVb&�M��ݪ`�����ߒ!�f�P����3nU~�
�����)� �5�����1�l�=㞈%�@���U�⬾�����Դ�:t���@�� lb$���g�Z�_2�i��Ftls@ 3b�~w�ɦ���w�c�/h8%	�>�cE�5z�Q � h1�H��I� t�-8!�+u�������2l�U)}4�d�$�O&�����)�i���X�{�4N�l���b��[ط[�o��66J�x72�(���s]DF�*U׾�I��}��J5#��I��<�0~�oώ���;��r��ى�m��㹕L�[	��D��o��_���������o&#�S�}��~��] �q,����)��[�l�I��� o	?���Bgp�8�?��0sg�} �Jr�Y�L���Q�����t��y���7Y�J�����W% �@
d{&c��
I?��	AJ�K�R����(�Ey���Q�3N��&$<5��!��_#_���l�=�heE���5�	Vk�pXkt�;>��Rc�]��;�E��Q�Y�k!qb��7��"mj@��7Ҽ�d�C+"�W�i>�o��ed^Ģ3-�w�v�V� Ck;��I
�%yb ��(]~��n�1�_�����T�[k�ː��j�8)n�/×�u���i%վ��˧�h��9�Ν����Z+|�e�\|Qk4�
K�H�\�N:�N��0z�L*��͛�ZA?�'M��ri>�3dƪi|��#D�I�7/d/~}�#���8���Ӫ�P��9�ʺ�'�f5-�����}���dІ��%��`�蠦5\��f=;�*��3�\M����ԃ���P�W��[���2?4ƕ�ۑ*��)�����_�v�)E|��������v|n���%d����Ԕ�c����g��!���>x��i���q�J�{,1����z��q�%��Zw�aglA�Il�w�-�%F����܅絷j�o�(�<�js �T�Z�|2�7�H�I�
��^1}#�\u*sId�?pOkn#�OՔֲ� 79�{
�������Ȕ�IC���TLmn�*д.<PY��{*�T�4���8˛��.3�7���,�x���}����N��Ԟ\���|%��Q�S�C��ό������
��| e!Л>����N�7�硪�*$q:�Aν@�_���U�R@��x*����X+��*ȭ�S��J�_�QN2Bs�	}U�8]Y;b<~K�)aX�aW�I�|1�H\F���Rla�Lr��C������M����$��j)��8Y���qR����ۤ#	lB=S0��I��YN�C���`M`G�_��Nu�l�D/�jt�;�( T2�y��wb���w����ޗ�q�~4%?�CQ���h�(�v��z�;ܚ,-�ʯ�[e��m�K�#5 �ud`��C��[��n�����%�'��m|�-*��R�cζ�SRl\��P"X�^/��=�S����Z��c�������f҅bK-��ip���2E+��A���8����ydZ#�=�}�3��N�n~�*�o$x����\?�AT�8DU3J7���N��{hYs���L$�� j����܉n��6�+c�a������������'Z��bݹ�{]��+MZ�NTR�bY$���aJt��7$�:U����cڤ������v$�j�����8�"�8f}��ԃ�$'�c�x�� ������WS]���Wz�V�r��ë��뱿�,2��=��`�hh�o�Ψ�f���;"��4H;	�xA���@(���D�ڕcA��ヅ��_�Ԥ�h/��f��h�lj�e�k^���א3�X��:���0 ��aHֽ�E��S�ƿ��B�^7�aE�4V��+Ƚ�:��DƋड©�҅��L�y��m7�+�����A�Os�༾a
Z�E���M�wi�r�"t������kep�P�rK!g�&���!bho0��A$�Ӥs:u�?H%mh�����n�1B�W�kP����=��p�x��C�e�g�]�s�KD�fJB�����y��,0q�WS��\�$$�s����d�Z锥>��B
��� &��ېW�z�5�׀z�.�m<���-0|,��*��@WcC}�F?�8p����Ҫ�Z�k�`��-�u�6���{�H<K���(����Չ�( ~)����'A�KZ?~���S�i^o���N^q�:_.���4�	�ie�Z�dț�`��M9&d���ȱ[gMM0끶��)}Y�/�9>R}��(�8�b1k� �u���<���\M�ik�b�� x��x5�~���c��q}ƃl���{t�� ����^�<3�o���)��>� ��͑-�d�}T��쟳ސ����n�T/���c��q��]����Z������tzM�>t�O1��[��c)o+�3��h׉���g������������*�ώ�j3�����K]��.��Uޞ�FF1���:�#Zi�����żkZ�LsR~�����:�*��~
G��9eFg�Qp�'���-!�6�/{�o*hj�Vm�ɲ�{;Hg~�:�_�z*�La�?A9|#$�?͛��hF��<Q�����t6ׂ�p�k4Չ_�y+�������� ���@���@)I~�+rTp��Uф4sf�Ds�>�޽��n}Y�"7���(��O���t�e9Fc��V��"\D���eMʢ�m�~R Q^hS/��k���l�R���Rxis!L�HF�BRE%P�°q}�F�`�\���2v������cɻE�A����|e듅=��.�W��9-�D(DL+�C6�k��0~E;�{�;�S3}:��;�*]��������j�ʍ7�𤠘ȵ,��9J�>��c����p����	3#���f�'ؘ�{A��t|^��W��	
�;�:�+���Ӟu> ��1�PY+��yk���$J�#YB�Z8ɓ�� ��ms=z���y��{�1�Y��s�U}���M=���hXr��_rU���J��H�o�x�ݥͨ������~�=�Ю��������~�3��/��IHD���]"�|��W�yc9+���~�}�-�����#A�Dd�5�扨�dUU�U>����-�a/�2R��?��#��81*rXFG4B'��1�vV�f�m��!\#h�h�	�k�މL�DȭD������v����\nOg�e9�����
Nٖ��8���]=�!��$����B�zڭ�+�-
5����yi�i�N��[2!�q�iX��9��W�>X�;�����{\�:u V�9�'_�^��_?�=}8[��v�2�3R>)����"�L'.i<�n�Y��w�茣o3�7�cH~�n��	6tE1U��� 4<�_��f��O�y�sŃ��+����~�:�INQʜ��-�K�X�JJ�|j��l!�U^��o�	}���qE#�ơX�N���5�����t���ftp�����L���4:^��<�q����t�X���rQ�=�A���z�>���J]�E�KNMʾ�$pw5�4�"|������g�uFl,�9�R���MZ����-���_�l��<���3�b�V:�ՠ������4�<���V̞�u�����UB@��Bf�s�"��v��7v)����4J���R�I\���Ԙz\*�d�a|ɏ�6B��QJ�fz�5ہ �Ӧ�<uZ����%���y����Oɀ�6��a��h����J����s�θ�Ҥ����=]��ؾ&IS��c�#Px����������>R#~$��r����R�<�xcߝ�ʅ`*���Fw�3vz�bW���
H���+?�� 7dB*.�$"�N�m�3D�aG��9Ү��T�V����_d�;R��+�`��J������Dө=�XM�"��A�����7ḭtn(�'M������)��Ta��Ñ��[�!����rb��Ӄ(1�S�'̖���{����o��~��h9>��9��'��t na_�>�t�0Zv=Ě4��d/Aӹ6�t�e;�r�jͽ�z����ؘ��{�u�J��j}�c�W�   �8�\�rs[�a�i�й-�A	�K"��S�s�Y�t�BD�#�ק�-R�'��7H��p�@33屿`	���t�o R�/��\��O�N�<�}�ӿ̈́�ɉ�w�D�%Z��h.�(�g��4�]���_��#�W����~M�0�[g.l(���=� ��5�0!�����c���n�]����G�~��BL�- SU�~n���/ң5R�4���9T��I$q0G[��<��i�@.�_N�U����cIYW��2�{����U~�J(��}�a�[�̒3;M�H�ើ#9
q����SL͟��W$H$3�؟ ���A&u�x��(���36�쪨ƸB}�ԠuQUZ�6)zz�����iUFD���[&<e��i~������<�o;x0����4ȕK����׌��z	<q-�E!4�<���R���VjIA�C������}�Su��K\�Q�e��_9��փ�V!���j��R�A�+(0��C�+ZS�G�$<]�P�EPIh�#�Jz�24�����EB���\�3;P�4�B�
ܛD��ԓ��(M���/OۓN�ua�����~�P}s1��;.ް*�S�+Rf�.z�F��/3�n��Ϳv������m�ܙ�.}����٣��m�h�:���Y��4/��痗�x�kN��i�T��f�X����Gg�G��N�Qت5��g��dN��.��:"ݖ��E�5��O���C=�����`	����l#s0i�wȥw�<ӝ	��\��I���P�sf!�LL:�	�m%ax�s�C*z:�"����ݑ�"-�]�_o�,*��#/l�`�"�7
���7޻1{ɪ~�,�!x�v1��b�/��7���J�t�:�s3*3�5x��!�����ʑcӯ�߹8��|ALؽ��VR��!�������u�M�'3�Dz[�J�2<b��ջN-�0_R����
llIeǍw�@�A����dK�������c3�1� Fq��h�&w��m����QO����#[0@짡!߾$c���F�F�"������Z�'s!l�C�`]�a�.��5z�`2�����i��Mm��QW`{��RV�@[�5������!���ݡ3�k|Mr���g��w�����>Q��3N�i���t���L���-������eP�y���|�̇ ��9�bߺ����C�ɱ�Jܑ�}��Ux�䕽8��#=�]8wh�ZA��H]�lq�"�^��ذ�?]k�.�ѷ��ܮ�p7�)�ux��Hv�F��n���Or��qY(<��!�tp�������^��«t|�lJ��r"�����k1.�#�����ZI��C�9bW�h���
I��E���liT����$d7CU�k{�)'K��/L��!��i���
�o����(�u�i �ٰ_�C�b
�P1�U�/�?�'��ٿ:��s�~����Eyt#��5�4�K��c9N,�c%�,���;ڽ�+)>��ǩ�O�A 
+���TaW��ks�T���E�SO7�]��ka�a�HҪ>��j�p{���s���2 z q#3S�5��-��X�t��q7�69-u��A�8C�.��F��޻̧�kW�J�& �p���Ʉ�ap�s��@�q�}�e� L~ؖ����vR��K���Rf����a{9��dƹ#����o�v���ǽ��A;z�	�D�$� ��Iq����$���9��%��UAn۷�s~Ri,���Sd�5b�����W�Cf]S����Db.E�d-QN��1?$�A�o��~���Lj��
��p�ab�	�p@�oW��>��S��.��R%�)P�j�cn
�����d�)OС��{�W��́��sπ����b����@5�t�����3��y(��8��9E�=�϶@�0a�]�`���)��[%���Z"��@5z�DG�*��#*{�}}��'�"��/)���d�N�U�n~��W���iN��F}t�y����*5V�C���P�t��Y_�l<>����4h�~�;�,XG<�n�D+�d��1u�Yp:rWR�1̤
/2hػכ(<�ɝW�p������-!n/����d�NiM�bc������"��V�����`�
D�|f��˾�:$D��iCPh��ɐ��>������tD1ct�\�N �
	h��@��A���Piu��PnX�,�����xAZw}^��jZ��4U�����.&�z�-~�O&��:]�za�1�ڟFA�	x��oZ���?U$%�����k����tSLF4]&�UY���M��m��]����G4<��*��T׀��ܬ\=n��M�2���>���V��O.�O�%B"J;�λ��bCQ?2��0OL�� ���*Ùyn��Q�&Z��/p�/�朔v�~����j�Y��Zs$c��h��4m�Y������=��N��o���fq�/~BAj�e<(8V+!��������-�4jT�5u��7�_���a]#zf�^��[�Hy�՜Q�v�R�{�E����|��y�l|�=o#t~���n��V�;�\ڈ:V�����2����}	���h��*��x+���z#��$qS?V'��)Q��]i���G֣)Q�17�K�G����(����0����~ajUv$�ie�/}�+9���Dz��P���w�%�No\��rנ�$_��������#B��J�L�}w�Q���(Ś�!��_�,R��_]r;���jVgz���`�$�O��+�J��\LG���b��O��MHr-�)�a{���x1��׸c��S�A�`�ۯ��y'Ĩ��0)���rm�>��~~�y�?�q�_��
^ʧ)">���A<�ׇ_,�>t�O��X~��w�q�6������L��l`m$���fS�7��?b��8=UYڑ�RH�u�.��d��S2T�Jc��<g����z��+�(�����`�P�İ��ǗE~6Xҕef��k䮔�k����ئ��|k���p�8:��F�(
~rZ�DF�#�������,ӯ�:B|M���']�dxDP#�#[o<p{�?�k�N_3��V������IՃPM��5,%>�Տ:�I�6n�}Q"-�G�@�λ��J�*'��8�2ڋЖ>������s�yW���.�x&G��ېُ֜g�Ʃ.cXؔ@��32g�C�=����������А;�ӊ(u:uP8 ������%yS*�z�n�������_m;��Z��0i�ʑ��xyk��%o6[%�_q4��&�0h���.j$=���-d���``�n�{c��R-z|�+�̣��x�ؚD����n�Ux��&���-0i�M��80�tX��N��8c^WvGOn�� ђ�F]�}s��{P�����q��S�(Gc׬}@{Av2�#���.U/9fN��t����c�װQ�Ԏ�zGgV��l��Z���5�:�H���qk+����/RX�S��6�qIN�B�����qRz��/Tb?0mV	�����v�ʔ��I��>�(^�;� ��G�CY��)�r���5
z�7�?_SZue�s$�Қ���2�
�d���"Ӯ/rt0��X+@Z%�����qG��W&Fs����\�#3"���*�vyЫh�_��2�Oa�u�����`��_�a�U&Q��-
��� ���U����{���I4�G@Ƹ��� [l�o�T�����zYV������o'�B��C�%������^B0����s?��G�-�UԗhբL� f"X_����45�S��κ�;�G]��=�&@	ݑ�E���[���e���-����a,��z��d�uƟY����m��09	G~s��M���BGӣr�ޙC J�f.�NM_�c�M[������*��;�-�Xŧ�;�v�9���ښ���!���կU����le��_M�߸p�N`��v��nR��`w���{�#�Aӌi{tv����8K�W�)��?,S���&l0��A�u?g��2��ն�ݿN��e�:w,qye�걃�Rs!4d�'3/�����܌)���-)y���~>���T9�e�+.%1+�ٶ?Ե/�s�CL�Zp'$x�����֚�9�����|CWQ��5�N���L�x����GH,A��<�$��������mO%�ֵ
偙X�ӂ�t��v����.U���0�vqz�O�r��^�F���.�!�3���8�҉�J�% >=_��u�e~()��Np�Q��ŭuA%�~�b0Q���s��<و%�tI"���rQ�?��S��x�,ͷ~�j�3Ra�Х٢�!��℡�x���9(��Ѩǧ&KiPp`7�=d��0�/E@%�GP��"�7�xϹ�%���~�|��J��ެ�8U���`��9/�2��+�϶���� 5̒.;�fڜ���[�¾?�?q�{.���q_��ѥ�{���	��6&T_�|�����\�k�?tIv�@wΡ�|Rn\���x���v��;��$4�M���Mb��(Yp�"�
߉�)pJ��GYRU��T0����ݤI߫*����;z(_L�v��t�`�
�"����q��v�뛐��M���L0'sJ�є;��S���4���;1�]�'-:��4 %N\wY������eL��4��V���^���H#t=e�i��^{�:^X�kA���^����o�._G��4����pu='4!
D>�P:.5���=s-@�L��e��y�.�7�1*�����+xpr�3g��t��B��BE���oT�����g�ٖ�~���ԾtO�>��[`����X��K�ݿ���9����8�1/3B�G��a�$���`�?�3wz��39y����Խs%X<$ Z�cu�p��E����NkK��ϝ��?���	��Lch�]쮌�~C�d��^��6M��:�ek0J�K�)v�O	�;o�6�v8l|���ƫ�e"�9��i�@v�!1�:��K��N��H1����.$�K'���0��Z�b&@W֑C��%�o4LNq�!~�Rx�7i��[(>a�I%i����l^T��iXb"����=(o��R��\�h8Ƞ �� b��e$+�*�]��RH�y��3��i�_��H��~�	$�.;B�K����ͽ%˙=�ʳ��TTۑYR7�s��~9N~��*)X�wCe���҂��_V6&<$nG�.��O$9[%Ort�n��ؓ��$I��]���?g��3NTl����ld�*�}��%шeM�t��2b9}3��0opJ��g~��	<��iu���h����^#BO��Z�[�����ì�9��TDԒ�
�Ҍ��(�?e����
�5a�n4�~����{������/�q{�V�KOo�t�r�b�cy��iM�\nS�?��k7/��ɫ�K��QQ⠉��le)=	��~u�I��U��>��+�bc��w?�Fn ����LU��pV�r��N��W����4��q��crMs��/���k�%R����M���n)=ϱY>�v)���ޔ&��1 ����7y��<�O����2�)fdt����'����tӆqy��
Y;=P(WJ7*������Z<B�)�׊!,�6�fֽ�X��h�Ē)���\�p��zC ����.=��A.�Л��z����|#rD��8���LA���(*��I|�I�d$�'iԸ�#k�Kd�w7"~���;@���&��/�쁝tc���P�b",W�\X��	>���K���L��~e��_z��;����V"�$cPJy�hxᣁ���C��g�,���+�̛)����y�NY��1A����ܫ�=�Z@M<���B���`�:O�m1fR�IR	���uKLJ�#�h��%�=�n���� ��
��k��p`����c U ��a��1ǋ 36�Zꃧ|���E��� 4�-�|@��� ���A�6�1���v���ֹӔ�W'�!G�Ŧc�A���J����N��g���{�՛*�m+���n�Ӂ�gEo�o�{�Y�o��������l�~�y�o�{	���K��#s���`4��`CV���b'��׹��_k~�Oᄞ/�iR�n�Z�$ż0[I�{rQ.l�DnzU|E� �(Od��<�Jk~��C��0"|q총��B	:<��IB���wz����y���ywIn[\=�_���j�����aX� ݪ'��O��Oʆ�6/0+�)��������mdf�������|V��3~`�H�bT4�Q`kw�ү�A�FK��}b�����Q/�5��ko'mq��n1�D�<^�R�l�4��Jq)��IQ���UMfgș(�8����1��J��;	?R��#�{��y?��\+�{i>5>�����4�*�Ц�x;_3^���W��Fb;=��n�Ks��G*��x!8j��d
����Z����ӓ��N̹��l��g�i �7����ޑ��H��N�:NJ��̞�opwה�M��ᮄ�������\ߗ|y,�){�j�t�1U�kl��!JS��
g�b6B��vh?a�N|݋f�w���p��c\�تhϚ�6ʪ�-oV���Fn3�ܷw҉v9:f!�£}�� ���{����|^�>d��x���՛7�6?��e�o��Ý���g0/">���=um�i>�#\|;�瓻�6�x����/S.�{�L��l�i�\T�\���'���wSD��}p*	�P��\����
Q��Wz�_E�`�*Ч��t����k?�w��ݵ�`�Z�S�&(~��㌂�����w����_�T��c"�뜎|&\���iUGUsv4TL��A3��
��R�8��b�&OV�.��\��^��0'
��# �b"k~~��Ik4tjV!�׍𣶕��C~r��?�-j���!���m�D�T���� �B���������c|��G�֭x+[���wX=��l>�9%R���T����Y�"�"�l���gթz��01d�T|d�×Y x=�v|	�� A�@��b�|9�3�l��_6��^p!]r�A-���<t�d�xZ҅p��5�z>۫
��%�^��H��.���	~}�uec�'~�}$�xInU埿�]��k��O��uㄓ8�b6��;�K����I��cB���i��C���^:�w��/��xv{�}�Ix��)�F����Y� M   G�m�LD�����J67�R(�<[q.Ųo�c�8��>r[C;b5���t��&��W�j���h�R���k�Ƥf�I�7�����{{n����Q9RrY�h]x�i��h�뗏]?4�� ��67]�%ԭ���i��;F�A��L��� s��|��$�X�N�9�?⣓1և$�h�!(�.FbC� �q�8�>�-"@_w@���(e;�D���12M�^<���� -��6�0öb;�1f�j��
}��A7�[��\�&8�񥸞}I	ܛg���v�c RKb�P�7J�ۇ81ċ�_n�Kd���B;eCiـ���8����}�7�k��~ij}���0D(t=Z�%藸ez�]Ԃ�
A+�X��!�]u2 ���}YH@�*�'w��f�k��EZ��� AD?hZ'�K[�+�$xd�d �V��|���p{�P4ۢ0��܃[�,zǧ]F	ː$��q�p��r�ǳ[�3e��c�����ș[B�:�n�s,�������夈���X�x��U񣥏,:�L��_ę����%�b膬?e��YR5������� R�3k�F���a���{r "~���GIb�BQ?vVN�yU��]�����j�"��
��eL.,a;/�*~
P47Hs�w>N��?E=;�ț�I�'�ˀT�%��_<� �����K�Wap����w@����%u����֡t��Wbx�Ζ@ܪ;4���0P��7p	$���}M�G=�����w�L�[���Ī�N*M��T8���������4��D�sPw�s7C/K�~ �����2^�"����7&90�_@� �ޖ���x���y6#C���(��N�<�Z�6Ʒ16y�JxCf�(j�Q��� �͝��u��ٴt�n�(Gc�0��r �R9�VC=����������2�G�`����~��5;���T+�``��i�u`�vKǉ�G���v��5`=�'%�a]�{\q���{����sR�Xf?�i�v��-�z@@,(��hվ�����w�%�@��x� �:�_�%�bv���γ�E��Y�؊%�~le~ÜV�p�,d�j��ē-4�W72��,�f�X6��x�u�'pj^����ա�l�ۣW�v��@`$Z��Ǩ�KhȌ�\Z8y��	�C|���X�Ƣ�hZ dSX1�tN�?�d� ���G#�����y����n~_�*d��8�ruH�:X%�A]�j�d��lP�֠����~��ؾ�57 m�i3%*S��m���+o���@9���6R�ґ��Z�Y9* _�]=��f[k&\��Vh�f��j﯐p��.)3WP^h�D��zK���C��{ZE�2���GV�8,Y�-t&e�B�������|�z��H���?_��Fʵ$z�f�fZb�N!0_Ow��Z�W7��.�������l6u�v�ݓԐ��ס� _=��/�Q]�l��9w�l���MeT�� ����~7�f��g��Ӭ�;��9�̛��;u�b��p���zF=�C�j<n�O2�����)�@U0�n���]�m����ݡU�mj�̰Opi�00�F]{�2��"XϺ���J_U��ٷr��uH��Ӝ(��������k��a�����M;J�ʠ})J�̮����*T�����C^㸳����#��`t)�e]9��&�"Y��Bj�3�ҳ���ّؖ��g����T��i�/�씯��:Զ���N�?�Õ)� X?8�7w Xb�*�Ę^�%��IJ9A��]���b�� P���$�4��_5gp�o/*���h�Ry|�� �=7�_Y���_�����[�ϟ�7z�H��`8�2�9��aা�B,����xwB:+\B��q�P-��a��=�HP����wM\(�T�9i��
e��o-�����&����q���J��nyd,�L���D���3�>@�q�ں��hֹ�g�(���y5�Wu����k���od�Q^"��:-�=#��į�	v��Mt[1���2����_��t��^0�c�w��jU�Y,>��k�	������J�Љn®gJfjV�<z����}}q�� #���͵H"�AT�q�W;�S�qHv�E�.���3j%3F���ü�RX�g�_"������gȻ�4��Ǟl�G��)�"�c�����@�x> @ؠ����SD��� Ƭ����p���tww#+z��D�l�+���B���'����	�`�:=`�����I�6����;�c��-Y��w�mr��)���0����`7�e���y&�K�EW��s�E;�ֻ{*$��q]��}G���hn��h�Fi�%9	��K|�q�?��c��4_�o���p��H���]\*�.(�Lt7����-H��\u�,�X�6{�'�3�Zm��/r�%�����q�Z�w5;Ԃ���wV,�*+��Cx�l�ga��I��,\lL��t�u0&��5X������L@c�f"uPFĉ�WR��7��xfH�3��E� �y������J���'�촼?M[��ki�Q�J<�خ�<|A�OS���\c�c�>g@�:S��E���q�=z�_\�?���3|�;όٔ��@Q9���M���4E���lL|����Y������ Ƹ�^ ��o����H1�(��<iZ���=������������z�
X�G�e��,� ���x�&4��R�"%�y1h��+�-5��g9ՙ��I���\:��V\����"���@�?�(���C���Ŝ��cX!��Ff�6z��F�5�:�V���(��H��A�O�d3X��Tg8h���lͤ�+3�
;��2b�6C�^��{��qW���N݆��@7����n�D!�:�
�[6�Z�����Ƀr�/�qɿ�]�B�AY��`�n��Ⱦ��qGy�C�!E۠{+~d��J��KJS�GL��0&��p1�ś��D_����ٷ��������\���'-1�]xqAX�1���-2��5�j������Jp�z�}���ֹ����E����2���	gY��Y�%������w�&����2�U[-#y2{���-���u	]��ߜ�Ov�=�Z"� �|��A�񸨯0s����R�X5���~��� �]���;5/�qYpk�(;()/{���׆w����eƂ��[#=����JHeht��5ޱ�V�����w�qN� k��S�L�py;)O�����~v-��䤝���.���m���⤾�6n �0��%c�	߃7���F�Z�V)1)owv"��R�~�dr�ṗmJ�t�x�f.����)v#!O�(G�0;v?~���T��^�[u��w����.FG����B�Ȉ�?[k���_���ɋ�v���o��P|Er+��x{�îN�	1=����.91�P{��!f�30�ob;���5�ٻ_1�4'Z����:�Q�Y�3�Xi����dt�/��۩��XDA��0��䖹��x�=6��)rnPB��Pq��fQ��6�zͰ�KT��9&y`�~5��^���g�>"���a��l5��͑��@��>c�n��1�,����(�K�����ݍ �O�5ze�t`���>|�y��Oy�p#3��='�o�Uh!�R➔g�$�6�ĺ��N��pzQ�x�����~Z�P�ח�؄*�%|��^����I���w;C�z�nc�����#}~��o(zZ!�uӜ�fMbF$��gZ������J�a��ٖSVB�b�n���lgbٝ�b�t6�C0�ЎЋ4�j���]E^`$��U.�},�f�D�����w����_���;�{���?[�} ��@+�<�M�y�9���4	c�M]l�Se;�kFf%I�>P��OU*�C���W��Z��B��u�&w1�Y���!��
*?��c;�4��h��կl����.����A�`x�[�k�U�"��U�T9q������lX�;3�G2��<Y1������el�KU��ú�ESޱ/WQw~�_�Д�Z���6W����<��E|O�ڃ����<lo�K�qA�5�r����e���4p�0����~JB�.�e��hu�,L~�Q�ֶ�V�U:&!Sa4�C߫y�Й6������Uv�ϗ��wN���a���G�b]������4;"�HEO���2<���\�����F��oL�hK�,�ig�q��0g5�h�R���]����?J�dBHW[�Y�SAMjY"��mҚ`:q��Q�����Zt՞ �_��}ٵI�z�Y��!t3��o�r���+F��ҝ:���a?��}�ǨV+HQd�&&�X3S��k� ~�_կ%g��ʒ�TS6�	�pK��i���]mf'��%~��
����<���C܌�EqC�.8$�z����`�]~:�ߵ�o�gh��J?L)Z4�[�u_Å�A�j� ��~B�gm�]~���}݅_��~Vʵ�KL��u��ME�����n2!	��eC.rˣL���*�DA��`�A^﷍E~>��%���N)�,��dL���������}�L�m��L�fz1�zw�v�a�w�B�0��=���
BSc/�ba9��j]EQ�.P8�8�Lt(�V<I��A#�z�9ԉ.<�����T�>��[D�n�b9��y�5p�3:K�r�::��_1uV�[~�����"T��0�|DmL$��u!��6�í������3�|�Wsl�[���ӱ�U�cA*��3b	�A,j��3#W�V���[��Iz�LRg��yw ��͘�]���|ז����k8J�d�h�-q۞��W];��TpT'2��� ��s���
9L�����%FI_�,�̓$~�ۙVq=׎�F4R�'����c�P�{��wD��NIWq�q%��'�t�i�\
ӛ�R~ؾ��AQ@m�qHS�!���Q��?��Z�A�j�Si���д����=(��~6 ��Io�+	#�em���rk9���Dߥz��r�&epf�ΰ�-&f�b�#���YCm��_�B]��:1�i|S�u��b��([A�N	�F-Z�H4���r��
��k��ҹn�;|j�PXBk��5-�Z~�SS���4���cC"T��3	�{:6k��M��N� х���׷��*Ka��O���ζ�@@3�2��*`a�$=Ǣs�d�G�i4ϴ�|V�t�S5*Qb��:B.#U����z�[�/�j��}��%��c���7M����p��#�;&�od*�c����� ي�=�y,}Ms<ŻUI�����h \q�E=�����?O�����_1����������6�QWn�fY�B{0��'�YXc9(�<�)~��%��n�_���/�v#D�^n^�Y��1�1i-����[����VÅ�2�[���k�T��<�?eS}���u)5ֽb)�O^�e�}�����1�k_X�Rj��g5��[�r��)!b[n��rŻr<����W1�W�]�zD^X�$�XG��J��	�5�8��bM���y��I#ENˤ��f��N�-���4}�qǚ�Kq
��N���j��>�o4^V�RTf��#���_R/Dk����sg
e,��9���GV'�?uBHH]u<�@���:��3+��h�|�aZlH���|�|< b� ���V*�8��|�'kz�]�D��R�Z�~S&�I]�z�����Px���tE3~����᨟�)h!Ʌ������\���?2��'�',5����K�8{��8��ʌЗ�g�vN8"�Pg@>Qڿ@x��� a+��"�S��`��q��Sz*�{�B�`����B����G��	YN�3X�s��k���U�Ο�����,�y�C���L6���4�QX�ތ�!��J)�椉/�q'sI��3p����n�Ƀ�7Q� �W���ƛ����°�1o�[IF���o��Q���'�y2R��RV~.��>r��7�'e?�/s* �(�z�y��>݆�54\Q, 8LԜsËu�@�o�c�!/���~�[}+!�}R�{b���y�pR��p��Ha֣+�6R�t�ҘCju��Þ'���u�m�,,=��],�1d%r�_�N�u7�L�=s���1vε��R�y�o�`��'��&0&q�o���I�<�1F���>Y�egɡ�V������_y�R#����NС���1�rj_7�U>4��s�{�7�u��5��:q1X�-Ln���%9
���%s�V������N����晇+���{��ăb�����/����P�-*B�����(���_���j�;�^��x�_|G������"��>J_��q��{jj�8�._/��+��3� ���������Z�$�R#� ��%���0��7S�E�*aK�sOY;4!)�y嶎x�%�	w�1ԭ�"�j�M��hmk�WDԢ~U�}��^����!�<̡"`_{�N�2�|�Gul��${������"�4/dZ�+29,2�����'�"+K�G���g�D�Co����N$�0V?�Vq��!IE�~/X[2>Ѹ��Ӿ�֐����C�/�!Z�,b�����s�/����3��P�H��bI3Di��|�����T_��`�\�Ϝ�&�����E���;�h�c%h�Y�&�t������|�z�Z�(L'�����Q%��f׆�6��H=�KIR^(�۔�w����I�7/Uv�Tǵ���W��[S	?\.p	��:���l��e8g��Aqo6��b0}�"��
=S���0��c�v���� �Z8�	Uں�A�!O��g,]�g�cvj�ӎ	'�9��R�6c�jH�M!8����Ug�g��@n�����f��� �.�p���8D���d*M@-nΜ�S�Hc��#)!�e�`������_'���cPyf���/\DC�Aˮ�3�`�uR~G��4z�W#�*x��XQ�؋���k���]�]3�癱@�>~�7j>4\p���ٯ��`Z��4,q9����آS(N� �ʛ��{�|��5�����5��y"2�7���7���y`J���2@�/�D��#N�ܝq���'ren!�y��3�{,��Z���`	����N&��?��U
�i�}�`�q�ź]�� Y���%��~���:\yM�P��6�Ĕ:���k���_��_쯲Ai�Rq�!�~:p�� �E"��	Nw8t�/�a�.M� �	v�"�&�N�jh��.�:Ѓ�c�x(�&�wŊG��J�G��#������V����\��Sii�OW�f�ST���Y�(��zlN?����^����<��͑�C��{�~�w_W!��ѣ�r�ڎ��膓z� �� mtZ4�����Qܭ��a�ƭ!��/	��T	
[	�`
ңT$Km��I;�)��G5��P=`0ҩT���D�ʚY@l�z�8�b�|����0n���:���X��3+��&�B�+�h�mu	G�-���6����}�^��Y�7.)bu/��4�%ޟ2>0�S�a�B�_�u�wo@�l�G:���M�oi�eAb���Q������r���2���N��9%��r)s%��˻�#��W���M�g�Q��$��~r/�:�aY�*�#��u�2�y�9�)��6@�J�n5�F�F_*z�C4}�y�_Wpv�~�<�fШ=v�w5��\b��C��q0φ�w�a��&�C�ߪp;��m�:���O��Q��m��(����У��^�zbE뗳!�ׄ�����z�Z.��6�[x��x�H��v�ۈ��4�ۯ0Ⳬ� H>w�Ј�)����+F��9 ���WP��{	�6^oq�)<���$C�t��u�j�
�іY8$^a�x�	�E�Q��?b�]X�@y4�����+���L ���. �p?-�e�9�V����1�e*�}���)�ׅ�!b��z�P�	'Ϙ��ٵ;�^�ǔ�W`
M��n]�hU�p�����y�ћ�,���TL9^`�@	���8�Cr���s�t'�M���#ŌLbOK��,�.��ROt��'}ѹ���}��LT[�/��f7�J�_�=?7����62�z#��'��5��bN����^����C��H<n�%�����dj�#@��?�Zp�U D�K�(c}KIR����7)��^�Y/�O�Dv����I��\��˼�/�7��R��A>B���_K����׿��� ��٣T�B���6-�IB�h⻺5����ېj��$��6��c�&6��׏cM4�����3�?IFp|z�2GA��Y�a���:`;��Hko|�s�ELڼ��d�FJ�Ս�\�T���X�K/Td_�
Ep'�'�aħ�l�w�3���p�I<���&��Ｏ}�K�<�)�a�Z�:;��?F����:RL�v%�q`��;��>��, 2Vŧb�CK�R�me�6��z���ݺZ�7������{�5��ߢ(*�b+��=[BH�fHO!=Ă�� �b�"��TEPTD���!J�
"�RE=���-/���e=e�$s�o�񍑕5c����BC �B'��H��a��Hh��"�[�Z�"ʦV
-j8�Kg�8[�@��xG$V�6ь�h#J�)��'D��:D �+��rE$�n5�X ��cY<��(��%a��p6(
)�0F�@�`�hZ%W:Y�j�1��h4"\Ov�:�"���F.� 0��:@�qz!��;!`�8\�Q������Ls�M�7I�X��L���H>0*�Y�92�P�i%���U��4�*�����hPLc��Na�k��H*	B���Xy@4="���QLo�tfI�p6�����h�Swci$�@�jԬ�� )�
����F*ĳ�a�����Qr�ʪ��:3Y#6c <3���j�(|#�,��p��#�*9YFrh" cd�i��=Ӂ0`��X�Jf	Y���dU˝.� �P�f��M�bY4M,�xJ2kP�M@$����8������VZ4*2���(*EN���@4Ύ
��تE� ���@��O�F�d	؆�ڐP*�6�f!
��pr��(�G#b��KG�" `��D3DDQ`R�%P���0"�v�3��\P �G2�
���p�0Q p�� 9F@� a�B��%4�8d�/�cX�Q�3�V��)�&��<I�# f��a�P�
/�dZ� )T��v9V��a�����Z�1J-��� ʨ焓i4K��Թp9���'(a��&`a�NV
9ZbT��`�B�|�T8��1P�Y�A�6.
&�1,@�KЩ�D :@G�� ;&K�
�D��@ 1,:�	k������@!�#�@��pI�Su��*
HN��a����`�s%D�4�Z��Ih-9\D��*	,�d"B$.jp�@S��E�
x�A�w�x�2@�������띞�a
I��lХ�"&Qa�MR ��2y$��N9v&��2#�l�)1�\��P�L����iA�Z�̢�w�U���i�@���J�*.ǥ�a6��i!%c ]� it�Y��t��;5d&��`��d�j�(��#��h1R��Tb9-ASH:���ċ��Q���@�O¹�( �%ȸ|�ZŌ֋�*S	���ε�sR�Jm����85	E�@Q(6"�S�A����D�L� 7��:ϩ��z����I8]8F��� 1��QH�(=��"�F�$P)�f1tr#��L}�^��@��H��vh�xAm���L��n%��� ����p�]m�rF�'�E0�\���@S�HV�U��`&7�*v���$�����d` ܮ�s�(��W�,�b��<�F�Dp�I0M<S��YH��T�Q,�-��vz���h����a�p�Õ�x��@32��$ӆGI�Z��!r�BiT$
��X���H���0����� ة0����'�l�	̎�G(�!� 7�U�Pcc�1��n���P�zXa5�lj�H�H0��á�&�@D"�jH �D�;��n�dD Xz� !��v�K` ",L��C�X8)�EPa R�� �("�o��QJ�ha�H1m��[�FAH"K���ŕi��C`w�9".U.��* �a#� x!C��@0,��v�~��a �j�Imj0Rm�Q�7R�,�RE��D�љ2^�4������-,1/nb;�0�N-ţ�%�pZ)D�H�Q��c����CB��Rf4��6�X�p�\
��D$��b�2�����P��#� *'������,�����PfK0N#�V��H�E�h���1-���Ӽ��6 ��1!9_�$Bb��Ee�\6U-��u� �F+���P�@.	�0;�:l -i�f�R#9�(C4,Ac:D4e51�4&��ĘL���XZ��c��9 -�����J�(WB��(G�Qi��`��ZE��e�@;���)�4

�Уqt*�@�
$Q��$a &�C�J�L�hE#A�z�>��G���%Bf�F�C�V��c�D��I��XRBB8�Kɣ��f	m�Ec"eF��%Y2��fW͐h.�EgX�|�Z+g�#�P1��d;D&-mBe|� ��IX3
���J���D�@"!� �"��P�6B8A�U�x�(^-0*�|9�(2�UzJ Nz��Er�,	6��k��(�FMR��6�Z�a��Pt�� 5v!@ ���2���C`B2��.-IF�(mBJMc��
�W��Q<A(�3�j5S���H:�D4�	2�X���)�
0aQB �d"��T�u0�"Bj$��R� ��՘H�1�(U�(5�d�p�8d@&J �k��XOa`�RU��W�	TX�#`�Xg�:���eXTV��.�Ѥ:�RI2(��9���k#"��@Z��i��	��)��@K) Q�H�3x"~4� 1�#�BHf�Gb6�)��t,!�!6�Y�7���Ѫ��\��" � ����S�"� w0�g3� %ӐP		���0K��2�Ёbr$���
#NB��p��&�[�%�(���,O�	�[�Q8��,P񅑑z��A���A%��w�"��H<����>��2F9�Z�A�@�8+d��B�j �$r�9H��C�he$S�b"q4Ӣ �ed��v��S����Ha�ɷ�M�E��eDj�N���2D��i`�Qb�V(�X�B+F!�,Q6��"�h�B��i޵B�����D3+B���"�z�D�A�(�L PA� �"�.�#E�Bd��g��� v4�3QaF5��$��RB��alv8��WE3�QD �S"�@���h,��"�I|J$7@aeI�2��ft�p+R�q��*�U��$�!��-0.�Ȧ�mJ��@h<;�!��$�X3�2�af�:PM��px�1�l�2�zU��N�2�5S��Gp)b!dw�QF�P�<�Ԇ ��b�	V[�61iPn$��0��Kdu�q|5W	� �TB�f��V�S�*=?R!dk�|��1�tQ8I�#�h���b�R���	t�"��w�M0���M<(%P&��lB;��ǈ"�2��e�*�
%���v2�Dar�h�.�j��b�C�#� �N�gQ�X���S�4�����h,��YT�=�n7E U D�ю  ���GcX:K���E2N�T�p�`D��� ,-�
��B��@��H"�(��:;܎'��Ō(J�s`��N�Rh��K�"�D0���Q4�N���!5t+C`���D.����l���uf=O���B0H�r��e�s j�C F�AL��Q�48(�lA�e`5��5�e4�F!���R$�-���T]F�r�mKuD�	� ���AA�HZ�1�,'KJg$`�@)J+���<ç;5�(d$H�7�$"��q�(G"��X8��U�-��.�p�"��C�y
R��:$|��8tb��J�1Õ��%�pp�ڦ�V. ��Ɂ�h�Գ�4����Ɍh0R�ߦd1KJ�X#��8\(�9h��IRH֐�E��'�h�Zl�6ʴ��V#��!����`�",<��ՠ�T���T�jE���dX'��T2$L%@��i �-$�1zy`��3�)Z%�ʲ���}Q��a�8�PCQ�� z�]�FE��S�j9�b9����\��c��P;�Q�8U�3کB��d5�=A��K9�(TFJ#Qx)����f	�Iձ�2��5aXFK�Mt����G�,:��b�t��R�dM�Y�T��n�8ͼ�a�<K�3`Y�h��;�n�B�D��� QN����x.�ǒ ��@%W�C��b�9�#��P�lxCe3kP6�&W��A O���lU�2� `Vͷ[$6���� �Zh��!�T)�8"`BK��Y�U΍��#��H�s��9Fe$b�Lf�B�I�6�̗�DX# ���,h:߆�6�ecQBC�ID��t.�=h[mS��b?���;��Nˋs5��e��������u���g�qcǏ;f�Xw7�q�'�O�4�}�D��ӧzL�6y�ĩ3�N�����5iʬ�3=gO�����MF�:_3f성c'xzL���ߎ�7]���6��:j���i�\���{���9α��'\��5�9�qn�'�Otv(��2z����1������lw3m�� Ը4��"�g��}'���_��E�}1X`�:�}��s�.Y�l���(�@�Fc�8<�Hb0Yl7�'�%R�\a4�-V�ݑ�m�����Jڟv���G����>��{�l޹�EW������߾s��������MϚ��hy����c{ǧ��=�}��?����k����;�?qMs�=f����p�m��ô1c��MG���������w�ҭ	~`�w/����Ő�Kz���?�����������jq��:ʙ<�i.a.?�슙~~$�̃����*{Jj��v��e����_��KZ�Q���4ʛ���+";�,��8���y98�����=�93P���t��{��� �����E�E��!7[��ny�ׅ4 �|*E�&���S�(�*z�~<A���`QW��#f	3+����)���N�^��k�k[�u��a���6&�������C���Bē���7�}�#���	����E%!���W�o��Yv(dE|�a�O��)mKx����y�)�	r@�s��,E�gdv��#�5�z���R�i�Ie{�Ku��J�z��\���׆���S�TPʙ,^h>��?�TyL����>¬�Cڔf#n����pv����_�^���*X��q,���#���LJϡϳK�� ���Ϗ^�"�>�\�kv��k�7�|n�_>n��궼](,d�G���j�[^_P>tO�:��Q�9n@L~�_��fL�c�UL�۳��Ԗ��n�eo�g=k,I�YT�|�������T�6�S{��Nz�Q��ȹ?Pk�I+I�S�_󯿡���b�m��Ț��)�vg��fY��7Xr�X�3T�֭�����Dxu��x����˼�qG��g�*�܅��N�E�ҿ�c.��_�]�.}�0f�*X�~�ܕ�^�`����Ŝ�)�V%|iɠg �o7�6mz�{g���]1�=�_�'�g+RN3�����i?������UT������e*�����KY1��v���I��@��=yL;�=����y������4�'�b�X�=)��u-�F\�~��-B���~8��ؘ�;f�v�Ev������W37����G�5����=�,���7;=m\N��~��ӑ���A��e^30</p��?���3���a��s�	�Cae�_%�WF"��hN%Eb�#���߿���K����َ�m���|�SU���>R�J������Y~w\�	�Z0,�{�T��@y��)�A�����Y�h5I��74��:�y�#$����vW�P��T�����]�g��E�r�aGqܝ߱�̟�#�n�����{��,�x��c߽���!��-}���m��ssmƣ�?��k��g,[�{�mӸ�jT�v�@��عu������d��u)y��벮�bu�R�C웃!���>#����Hfp����P���ۑA�oyh���OY�����?���%�F�����A�թ7H��Ϣ��ֹ�=��W w��,Mx\-���S�
�oV���y�����to{�v�|�A}�2�g�\�8ݷ}}��-u�uoE������ہ����}���.��~܏� S�����0�/����?r��X��k���_}9/�u���+��zt�����<�7��pS\Wr�&�7�lH'��a������Ы?�W]��6�fQch��09e���h�	�9U��_�Z54�g����_�W���?�o�\[�5L�������������#�d�ظ3er��g�+�������q��-|Coa�(��LY�����as�y���E����{ߎ��^Y�_ڴ���$�����L��H���ƁC���k��c%��m?W?q����E���!O���~:!:E���oߑ=�]d�!��龤��9>F!3
#��j�����)�O�ݺ��0e�N֚HG#�y~W�w�ι��W�Q�m:�x}�bur�{�I��]����l3G����� �L?\{���`Y�w*�cd��8���� ]��p˯��D�ϯ/�K����ܻ����.W��_O����ZSW�p��;{��K&G|�b���c�<J��!C�S24��yg�ג����㻫V]���C���2֓��o߅d/����D��ʯS]S_y+�֡��t�m��c��!U��m�v6q�m����^��	�?�%~�������?k�R[�BdW�������ʖ�\@n+,͜<�]\sk��ђ5-�����͠��9���\Z:�@@��#�Ň]e~�#��_��o�T��L�"�4 ��Tm���K��������e�P��tYq9�ρ�]	+}dU��&�Tmp��/�@}��iܲ��g-�v�n%���;g#/4ߩ���yu��64}�ԟ:Q�rtv�w�5�{f1U�hRG�$��S:�7�x���-�H�)�R$����?W����%��c7�~_��и*��>E����ߕ��	������;�׆�wz����
���Q��* מ�XB�'�J��.nL�1ŷ%�������g��I��^$t�2=�q�>��������g�w_i�61�<e̚W;:^5�����+6��������P�+1/�S4|��7}%R����_0&]���A����淮*M���o�]题Q��B��d�L{Ь����gϤ�?�1%��B���}�*<���R���R/�����7�������\G���$��y�|�Ş/��%w��"�����yds����u��`�����\㾡c��Wi�̒s[?�Sߧ�.s��qi�	?��qf��V�����y������{RΝ`�O�����;�Z�׵�r�\|' T�~yJ|=6�{Ҙ�ޯ�<����4⯊�w��)��҅7��X�D)��퇪�����7��^�����;�_�j��p��M��ϛ���a�����ӂN-�r��g�ݝ�xn�W�b�A{���X������;j���Qw$�˛O�BW���^�Е�`u8匚�o�f��7�Pw�.5�jg�����]��5�n?��>|��񓼦n}�b�Hߚ���o���y~����n@���� aO����e��U{�9�&�:�Hٵ�{1f���_�ō�O�?��!
�O8��h���;n=^�_�u�eQc�~H׋���k�\�o���_����hwV��g�b ��g��-���E�&�=p�1�����%G����|�<���d̻�c�y7@�����Ԟ��6OO~��u�y(�x����kjx�v�b�uŘs�ئ+�t��4������17�����(�H�
�^�����7;��z͂��g��_z�V��f�#��m��-^�t�Ėʙ�q�I��w��Ν���;��Rl��u�Ԋ�����x��q��"~��y;�~��� ��{�~XUB��ԵNr�[t|K��q�CW;ߗlD�Vn�i�7�ɍ�ڠ�IE=���]V��Yh�j4ʏ�=w��~?g oVu����8L�mڜ�gS��w�m�ʍ���_�O���?�������>�¥�������iE�c&��<�4BH�[1�5tL?�8�߾�E'�6Ο��Y]&lS&#\�b������ץ�.�x����Kf��P~���C�i��0���zƞ��qCWRSbR�c�U+�mY8�پ�K]^]�ߞ��L;k�]?�{<��_����3��a�������u�jhG���0{T*O�S����Cv�����x�Ȫ��}�.j���?�ɓ�g���:++����J��|��eb��Ą�x޺�C��u���r�7eř����o*��G:&���4�]��,��~�/�����.?济q/�1Z��}hWP��Hjܓ���w�9�j�ů�1mA�ĥA4�g�_��⪸���N��0q�\��ώ�\���`Qo�~���e����=�*���7��q�p#���jѲ�3�0Ij��VV�ی�]*"��l?�����9NQ&�`����;�� �x���Aߵ%U��EJ|��NI�{6�rN耳'����|׮���I+z��ڬ����ZP2��
~�&��s����Xwg���)�{�0Z1O�<�s>�u+ص�O񣘸9xt��)𤥪�c��r�닄_���U����O���v�b��x����ׇ�Y/A�>�7�&���U�)������w�U��L�T�M�1-i+ߙ�H�eY�C~��߬�u<�<�}}��O$��m;gJ�m�+Ie�P����4}}
��j�D:rzw���.k�H�3뤙�S�����C+��U���Y�FhdC˪��f�H�{u��_�������}�M
j¥/�'�N����O��i�1���|�+�z/}���rȵzo���/�Ŝ�����<ͥ�y�_�_M���� ��+�|0T:O�3�fȁ�NrmlM��y����+��A��kf�� {^m�RU�U^��e�@��:_��Ǚ��I�(2�v��g��ꯎ�c]�o�W��ƶ|0�����u������A�~��lI��7��u��{�c]!`���\7c��[�	�NlO���������FuЎ��L}�?��3g�����!��w-������k=�]K6������Я�s5��]��3~��KA��[;+�ASOw�>��1�.�֜(�a��t���ٷ��u�$Ny�w��L݄͏��3{]�\?�v{熢�?6�^N���ԑz�M��_b�VN��x�gjy̗����H}	I�Q%_B��F�I�<���@&�:������RPg���O�}���~�=]1��������{!]�ac���d,����3����<I8��++cK}yK*��\�(L:9���9�
U��O[�dM�g
3����]��&7iH}?�i⑿.q/��j`�<��kZ�������Q��P'���v���t���/�?O%���!������0�"a5!f��p��^��=*B����E�=������6��0���.��F
�ު.^� �J`I�עv�y�����
}�3X��ҟ=���:�سD]T�os^.f=V��s��g\X<�����Cc�J��ğ��rn��U�Z3.�<
P���s�-������f[���is�F�j��or��9.�/�h;�y��hQcC\�����/���}]n��+�+M
���K�ph%�4�R�� ����r��8�-j����V1%G�1��P��ZH�\صx�6�9'�U�MK��͝{�ǌZ����Y�����T׽�H͉J��aK#���ݩ.���T����5--�i0�N��/��˟��{�n}Y�u�R6tI[.�j�o�������¬8���p�[XUR���E�Y�)j���ܳa��m[�*8e����������՗f�
�5K���+��������5�w�	\�����C���$���s5��6�V����ze�����͏]Z��xU�P!�ؠp����&&-�3����l��������}�-ns {Ύ�Yh+�����)E�M�w�$����@�:5���8�x���'^^��C�cm�3��f�Nm�@�2^�C)��2v���!��>��C�;r勻;jM>��;����@\�Ӗ���Y�_x>A��~�\�29l��Үߜq������VÔ�� �G��7���J#4֩��+2�=��>��c�0�٦����m�_��o�)��+|u�Ћib�y�ȫ)���z�4�g��v�IO����-:X#���IX�9Y��1��V���M������~뎶{K��)�z���}���?��W=Iy0�*\��䷍��"������le��_���0�j�����&�]G���y��8��9����+��z��2���6�	bnw}[A\��0��v�R:���1k�H�����9�4��c���Λ����z�{rC׹ .�i��܃��:Zn���q���]JFsÆ	��3����Ⴂ�u�z�ܽ)���们����IW��h;y����||���S���h�ў����3�Ps�^�D��~�_P�m�U&���"l���\<��'�j�n@ׇ��H�<��~��p9jp�����o���S6g���+Ҽ��^���O��>��z��"�i$;�by��=]�Һ�ڕ^�O7�7aɣ�<e��[1)��͑����D��x]���_�Eٖ���^k?B2�ꞥsܒ�a;σRR�̧��)�믧�Xݐ�"��6y��͕Q�Y@��4�x+���c�I~�AD�m��[\�f�Y�mY�
ȩ��'������Μ6DRc8�����S���N�[���Z~d��.z��lU�b�hKW��+3>4=�Hʇ!�M����ggү���Fb�u��z�������#Y���%QG
�?;�&������b[��6�E������gkE{ۏ�"�d@u7�q_-c'ǭy^ r$����y�*��8_n��g�/Ϛ��E��w�f����M��Ywb��*6xn��K����\o��A�9�wf��J��3�)�e�`Nkh
��5�g�qKb
��3�`�̷mC^k�<�gK���z5mI'��y6�/�Gi=&k�}aB����u����8Pz��"@�~*�e�J��Y�����L_E_�m�a/��n�~��y?��;��x�|+{�^�J��φϡ	s|m�o�4�r��ĮJa��#'q�WW6ܘ�"�#N|��_��\�O�?���t@��i��o����G�װے~^���/�x�1�3����̬u͍Y���^���oa�G�7:J=^�hW?S�9��BnTʑS�27E(j6Ik�VVF��c�z��~��T������T	0�~]R�t߮�`�`�i͊��_�C.��y�0���5��5������YhZ�K������_��Ȱjѵ���Ts�H`S�l�{7�l�n/=�?�~U,g�*�r�;x{��Z�{���k��o=fZCd1oF����%_ГY]���G,�������㵋��Z�j���/}���}�h����K=��}��g�� ۊ�Sv�(�;t�����2�P����v�h!�_�qx/�}K���F����h�"�_��:�!&�ր>7��l��mKnhM�`L>د���'��0��҅/��[��d���^��\�ф�Kpx]Rw������~��\w�������&bщ}ɛ�s�����/~wi��n?��{lc�y���b���9uC��r�$^&~c,{}�
O����2P9���1�{B�'w��<�4���U�ݣQU�V�(�ʢ<B��4*�mFu�6.�{�D��s�<��0r�N��ij�c9��G�������z7V�/&�Q/�R����8yT�,j�y��q奘Iw�����ڵ-��7��Z�**m�Sۗ��!��d��>̅�x��zm��v?K6z[�:y�n�@���r��e�&V�����s��-N�Y9�Y��a��UGr�Լb�;ۢ[�I?8:i��K���eƤ$�u�>��ȹ�%F0�\5(�˩�r���j����u�̐���E_w���.�������e����bvͼ� ��l�,�����>���4�p"����Ǯŕ�{�U�ꙙ����sn!�S���<�?rI�^�ӾF.��6D�.*ϬZbx|�^^1AXR䜏F9��K�?m�����='��zzrK�k�y��h~���<{��b�{p�ڸv�:1>�^�!�ͫ���
[����8�����a��B�Э�ӎm9���}z~��rkғ���ޥ�R�u2w���S�׆�<Y{�p�U��1Za)��o��\��|R�\�m��#0�:𣏕��-���B��ކOA ��Oެ�~��"�/$~=~��m���0ݷͽn|r���שA�k'[�]阯 �G�$"}��QAf}MNo��-������e�sWk^W�р?d�GW��_���-w��X���k��&�T���{��%i8��]��MYo�����G�*j븿.�>�����=������~>|+$3Vȓ��+~�f� C�׮ͭ-���ڑ4���z�ɛ�c�C3����㿎���Ѽ/��U�/O�c�X�|i���|ֽ���8y�@�kes����)n��{�*gR����+���7�E�!���W�g=��¡[Wo_�|��)��ܞ;�
B�K��m�s�Fn+�e+*�h�:������T���-�c�P���r�B��o1[��WS��K�߸� t���W���;����[N���^p�ѵ+�u�#�˳a�mnw�}�;�59�S��qZ9弭0u*ٻ��G�qn��b��|�`>8��x#��<-��$������\Ɏr�Z�S����g<�1f*/�g=|�I�+��~zT�:���p�:�{D˝EU��i]��'�/��ӫ��ܦ���3��~8��q׆�¤�S���}�oK���l�Z:1VR�r��g�[��ҟzu�g����L�n܈��Z��b�%<+o�G�����/�\�Op��x�-=�z���0���`��c?|Cq3�Ծ����㝚�8��J[�վ��R�<����}�t���t��ru�!X�rwYp;��_�5i99ǣ���>*Mn�f����z�5P�΂�[J^>���0��+}mg}>��ƃ�O�ɂ�0�2�;J�W��+���R�L��iw��-aJY�BjN���io\j��y֙[7'�~����ϻg��>�ק�>���:B�4x�j��Ϙ�݋3AI������"?���h��q��*8O�A��b=4;��r�W5�(��ק�����w^����ٖ�9'.��Oh��?W��ّ9P=f��"�?�=���~��^kNz�	���b��")�E�e�����R����ӽk;iF��*G2�cκz��8����ޯ�ZOK��+JH��7��ۋ�Ӈ}ߟ���F4?�1���ga�i'�bR��R��m�K��nwZc��xA,A��>�P��u��lz��	pvH��&�ħ��$�N��i����ЊJ/~;^�{}���>S*�~�$�њ�����π4��;�
�8���uq����ߒ~Z�u�_9���bP�gy�����r.�~�}��[]R����Q��7�v�}4��A����^��EJضgO��M��&�t���!j?+�DÁ^=ఖ������m�����_ߔ:���tX�*�[�We����u�	�/��{��r����K��;mHɮ�ڰ������S<hF3{�?_�9\"��P�CZ������!��Z�u�N��8��B|������M����z��̹�y�3��4g�����M<�;����B���xa{���OQ��7rj	1�f�%��X[a����.{��/<��E��V��ø�C�5�<�����9V:���}}&�5g*W�u�ԯ�6�>�e��0i����%��$@��ܵ�{7-X_���!s�-�r~hW�2��_�i���U�'ǔ����<s��f\m'�!8Z�b�;7I��.��@v0a�5�&�g�nxf��hE�:}�s5�I��������֊��W�^����j+��7Y��rN��U�1������5��KW]����)4w*�������������u%���'����>��6���Qޓ��>��kyz�c!s�������� �1��;�����Cx�f/Ć�9ˍ��S_�R����N%��|k��n�.�K��yo�[�c�T�_.���p,�,�c�<�
{b���޸�s�V�|I,2��Ы��W=�$߲�4�����B{��w�y7CkS��ܱ�Kޤ$��ҋ��Ƕ�?�z©�ޒ��#۶$��H�~��S�V�߾g���\
/�#��sM�7�=�r�`]���?Т�iSA�%�,�c[����\7	�>�w�̾{ˆʼZl�[6�sB��W�{�$�y")����s�4y�H�w��x,�8����ݻ��>Y9"��9�-�?m	����Z���9X���H�ݽ�챇q�|�\|}V@
���PZl�?�8[��^]��X=kiy��mۋ��O����t�r~kM�Vu95͵���?kJ����S�Ĺ�U ��O
QL-�$�� 
�v��:��TZ�FGģɄ��hz�-A��Z-]}��s]����:1��� ��l�����vK!�2CW�3`�~Om�=��kݳ�L�׬��DQk�ʁ;� W��F�H�V��:)�ߟU��p�{d	N����aJz�En�{�0�Ѵ�^5h���#��}�>P����+�hL��|��'�ܡ��=x�K��'��x��_�g80D������=��� f�<�:
���T9�[��pҢK�?���LD�:�L�<�l�2��U�?�&��	J�ۏ��5�#���g�@*	/�݄9C��Sޏjn����'}&�=ft�����o1��Y�#7)�������/��7�Y���g����N�/	�� l{xu�r�3������'��;��~}R^�<�����	�����}�y�V�'�i�W�w��a�qNR�s?��R��l�G�p:��n��7��9ԑ������՗5f�xǌ��%gyx��]�i_����)K4�^�Z�i���Qa9&���c���|y���Xr�	�`tRs���&��Y�a��2k���=Qk���?U�t�d]������	����J���������aω!���nո5u�����eS�	ʳ{����[,Lz�}ϞT��S�lOz^z��Tnk*�ĩ�e4@�G�ǅ?2��R���/�ᡄCMu�L	/�~ʛ$FO�X�3>	'�|Z�G�+۝��Dw;�P[ʕþSW�f*�[W@��))�1A�P6�f�yJl�����sz_nڥ���R�sCtt��-��_���J�^Mr�����K�,ٺ�_�_�$�^�v��ռ���P�NZq��OJ��ދ~�//k]�p]J��k�w��>RW�o
mS���M�CIg��qc�1��V�i)W@�f�n�F	0W�N���o�� s>�d��������U�{��' 4ǿ����^���T�m۽�7S_��{u������f\�G%��R�����'S�3����jm�n�>i�[�>ɸ%f�Hؐ|L=f��u>H��|�����9���%��ޖlB���y�uٷ�A萯�⎙5/���C���>�Ԅ��n�;
�1�V��)Ѝj��}�H#��f�-t��r��.5�8�6IuȮ�x�����-���e{�Z��T�!���1���������v�Xv���.�f��B߇5Y�P�G&��}k+;8qגR��N�̇�i��x�)M�)	������\����̧s�[�Y�.�qO�ϟ��L��[���T���o��F��ce����'{i��'%���P��v���d�}�>n3�x��z���G����3�¬Ы���w72a-���Vn�W�J���PSz>(��aPO�a΂��9Cq��w�Q���m]w�ؒuFޱ�-���:A�8���>~�T���4e�y�*�w[z�O�cq�8�;�f�d֮1������O�\�劘��O햡���A��I���ENL'���蛔�^����撼�������B/��cAHj���,&���4��s��?�K����kܒ,�۟A�`⇚=��8]��P��K�%��J���ΙN�]U6߃ɽ݋�>+k3�D�ՙj\��13K5�ϓmW�T���vոɊ����y(�<���F���k-}}ov���!.�w61��Ӷ�?�@�r ��=K�X�]�I�Ȅ�z�'	���/�gL%'=*M}<P��s�[R��eĊ�Z�7��f���x�;���J��� Ms	��Ɩ�à��i~��o� R�:��,J|x�#�A'A��۸����zζ���^�MV0r}�ϖza!�;��	�h�x��}���,�>��7�ʹl}3��(m������ɵ��ˈ]��Gq���m#����Ν�R��^��a�1i8���S�1�˘�������_0Էn�乗��	�_=��TQ"�����=v��������W4��OjJ�:L���YA1�� y���_ �R��?��6��t��ZK�
���3�'�Y����E{Y�X�~�����c���ٖ٧��c��?@�����S7��9�<H��`��iʡ�3�4�����}��1[���`v����L���� ��=q_7���W��ډ�� W/�g~�>��Q����Wu�}(��g�-��� 7��܀q����ۖ�x�J����MR?w�}u?�)W�dM�qQ�=�1Q��M����!89�:��j�Q����BI�g�T=�BR��P�i=X�OʤV��LU�)�C.4u�d֣��+�?��\=����G��]bu&���A�m�{s�^7s���(�M*��k�@�/i�,Lp:W����A����0�I#p��osՄQ�V7b����+���
֢ۘ�׉Y�e�B�׬|;�����6�j#&m$z���OC��^�|��#�+��B���3C!Wsf~�ŗ<ӡ�.8�� ��f=�kN�IU^ ��*�.������w�G�RET:-�y�p:�u��2�UEf7�#^P݌⣺�Z�����-��q���WR��v Ȓh��ۊ�@�~�EY�,�o5q��T8�*�?4e�Tn-]��?
��Ñ=�^���k��Gb�rF+B�ܨ<t�]7�?�^*��2*?,T��k,��ִFb�&���T�d�1LWEFnh�{Ү�������)�R�\���:U;�y .A��m]�~�eu<�
,8���Fq�U��$\���+����9�L:^x����q��{�A�H�09�]"骫�9����G4�Esl�Hc�����{g `R}��'��1�������-��q]�v�**_����r�nymǄݟz�I|dʘ���z�����1}h�A�����!s�To�#����8*	-�E�A�������� �=+��� ��]��Z�ʍtv����n!ڣp��N�,>�g���Ҹ�h"=�nn+����Fk��Ԃ8܊mh$��%��̨9��\��&�� �,�3��k!Qd���ԫ�1��^� �5�q�Z�m����k�H	x��)lz����$玕���W�2s^�o&���x�K[�w#>էC#��̗j��g�{_����1 ��b��t-�rq�u�ahYT
F��������|W�� ~U��&����}��q_8�j9k���K񣎮��4o��Iۚ�]� �WA�|� lHA�*��ͽE}����O�37|��{P��SX�k[����s�4�m�R�����zRx�M��jH�zs@���nc�Gj@�恎��9P��tl�,�@d��џ��d��k�7ǖO����g�A�~GҸ1��`�#�KbM�J)m��<�Q_6֧ѭ��//�O���Yn9V�������q������p+��+W�ewa���FiY�
JC[��%9��Ҡ�5�m3��O��piF��>��!��g��)����9�E<����{T*�OLӄ�{��t^b��d㖯��έ
H�5�߃�ۭE�2��������#�+��j����0���붸�w�J��u���A�+��$<����v9�]4It1�5��� �\��)��5��y�d��Kb�t�|���L�U�8滻���q^y���X"�R��7��c޶�i�e�\%����Fqچ��d��O���\��4�ul+��A���k�<;�_G"����t�L�����UA�E
Bh��Aa�z
�$���_���w�>�i$��q�W�W_Uf�D�}��]
73zhi�Ο.��}2+Mu�.�jc�5�n������	�n��� �Ԩ�����5W�ϰ����� ����9|A��Nng���|pE�n���2�u�)��� ��Tخϴ��(������S'�,$_�do�M|IǈY��G^�x�e�&����᩺m�2����r�?*o�$�K��u���� �L�cޣ��2���A��8ػ[���Z���˻������W���Q��#�+g�S���[�2���[�V7���?�nCKϭB�$$v'"���b/���Ċ=�6��e�����-�e���c�<TR�X����֜��>�?, ��?�ޚ�,�� ?�|^~+O��N=�$��3tv���_3���lˀ�F>#�s�Z���)\6>r?�O�WH�٧�.T}�� *�[��j9�*Z���A��3� ��u�~v�޳u��7e2�Î��_A4��-���#��W��^$\�k�=k�U�3�\������ X��k��w#��R|f��z�β/�5,[��pگ�� �u^�����j	>,_^�<���5>��A�#�;���0}�}3��U_?����������j�����K�JI�~��Gō
3I�֗Ʒ?h�bj��^#�U�c����2i�R�V#*ErK{����Oot��3T,5y
����Ms�0�;?�eC�����s�7�V8�K=���{��X�j`���U�����8�B�t!�#��2d���ь�;f��_t�洢�"�N+/R���L������sM�o1sT���5kJ���#{�o�lzW��_���_CZ0�3����f\q�ס���Z�
��� �o.=Ms���G�۫I�>j�ZLW���Q����w�R�cMFd��� bx�Z�ْT��Uu����R��i�v�#�V����-Rq�M��)i=0*�y�hq�qOE��R�Ӛ�C%l�+��h����Z�����d�� L����^�;�zH���O�D�UkRV�6>�W�D�?%�Q�x����[�j��YO#�N�ş&�>y�����M}d>|�o���m2����#/ҙ(m3ni�I�5%!��~��ny���4���jM�#q���t�waHƳf�
T�i����{R�=)���*F��mZ��;W�?	wl� ����~bu�A��b���G�m�6����ᗸ}%�i��h��_h��3]07�z�V�y��֧ׄ��8#��oz�{ć` �\�B�&��GZӳ��$q��,���^��W�j\g���M��H�\w�]%����v���	��'c����+cg��*1��yxJ�#��\��Ho���>��E�r�~풵oR�T��v�w��m���'�5�U�e�t�56|��?>�u��=k��%��(V9�����}Z�ѶN|e⏛Q������Iw1�v2!�.#坾�5$��ϖ�����L�ɏ�=k��XÙ�ou[�$�Y�A�K�����Iz��j���4�P��j�����l���Ez>�p���LדZ6˄>���M������Sw;vf(�cKۮ}*��E�d�6��s�\���d��7���i�?�U�dm������*�ڿZ\��dۛ���.�=�T�R�GQ�W�oQ���O;-�O���Fj��)�� ֠�>�W'�s��;��m���D'�O툱�4����ZR� j�z�rt4�j
�Qs2�1nk3X}���_$$���Yzֽ�H5Q���Ē�8�R�ֆ�x.�����#�o�d*��5�j���֩���j��H��(H.ͨv�8�67�Q�Q�p�-J� r*V�	�#�y�-�c's�o�����������:VK5R{W��|Y������3�_S�P_
�y��:�s�M�Ln��K�Z��yz�R�y2Ώ�Z�̃���S�	��*�j�S^H�!PO��L�y>.F�>p�Щ��`yrβ5RH	��/� ���s(#�P��Bne�Ӑ^�qpU[�Ig�6 ��_�v�r$R~�j��=����9���Ȟt{����������>��G�5�fW����\N$pG<^�����Z�V>b��� !g�L�-��nx��o�){��n����>^����P��L�+u�haaW�?�Kۚb��J��%�/&�����c��!�=*E�S�nM=W�`��s�}iѷ�3�>?j	d�yK�WП�['���?8��_ ��k�d5#T����~�Ŋ��/�}�ol��b�%�g�Q_:}"Z�. ����c��!������� �����������0;�r�oZl�#Szv��n��� AhO4/�E#��۾i��K5CG��MoPiO�L8��+l���3�L�y��NOzL�f��dH���������ǍR� �03_Gp��Nƻ_�@�Md�õr֧�wR��~�X�NI4���(�k'T����R"�;��L�������n>3O)8l����ܫ.��w���n	�+��L�H�s��v��.�+\L�+��Mg��"�U�ȀF5U��=�O�-�&������ �]���Q@�G���$��s\����$\�B�O�4}ZA�϶���c�����>.�1���U���W�=����v��y��cƥ�h�QoI�soI���uϊ�2��v���o�߱͟ƫM�
�^<���{s]z��ď�B�dݞ:׌jש|���8�V�ķ7D�|��r�I&�y=MtFFNwЛ��H�I4g��ӡǙ��т�8d���T�1FE�5��s!�����H�;Nk[L��p{���@�x��`�rMZ��j�0�5�r9�2x��Xw=M՚� 9�wWL�3XZ�]���MJ`mNO�Q��x��v�Z�o7bqT�ly��˪ؓrOLѦ3��sG�$��k�w�#k�I}I�-?Zy��q���V������AI�ŝ��`����㌷�3G#g<�����Ȩ��z���Ȳ~H�ˍZi�i'��X�=*�U��<�i8��t��	m��w�_��`��ڂ\����M���20��W�����Ȫz^��$�{ջ��=�{��ZѼp�L�b@ϭz��d*�z�ׂ�n�c���kv#vE'��Sq>�� ���/���B��|����_?ǯ��L�%ea�/e�f{��B����:��2�~�7>��v�)���#��ժ)���,�A<���<�������!z׀A㦋ws�Z�� ����ֱ�ݘK�{ռC��r}�J�R9Ff�k��⃰�r�/�-��a������=��}7y������{z��� <V���brH�j����B���@>���^=��ٳ]Tp��Sua$����95s�/��;W��C��݊�$c�5�R/ݠLT\5Hi�Ӎl�Q��I�
 i��Sמ���R���T�r��չ�~��֚'f2����եS�?�x3`G�^��(f]Zpz����_ۅ���t�6��L
)-P��~�W�=ϣ�����v� �s��f� �VǎT/��a��Xr6�N1�������9wJ��Iӽ1�*l��IѳN�ҤЍ�f��z��j)3�=�6m�L�������ۆ�y�jcz���5AI�g�����H֬L� >�.8����JX��j�`%�J$�zf�ΐ��jX���I��ӜqI��F�;�i��[�}�U2lbNsR��8���ۯ=+�m'b��j7��"��t{�TMʒ;W�:���ri�a�Vm���g�ޠ����k��!n3��[��z�}���=G\zRG�Z��EYI���������#��DɄ���(���ہⱜ�����9n�����<�r�#��N�i(�b�w{ֵ�3`�9��k�t@2I���ò�k�0��McӠ��1 X�j�g�Τt5b�=��rݪ��#�/�NF�X�����Bҷ\Wu�3&1���2"�^���]����T3�Z�1�ꆛ��q�J��IkTVd(O$qK���\�!��Ԥ��>�),c��ۊkD�W�
���Ժ�=�7PV�Y��@q�Y��~ ���8�c?/ן:퐮9S}̆��=�@�qO��zRwE�{��A�ռ�f��\/�����ԛ�	�]o�-�k| PU�WO.��Y�b�����1�W��\���M�)\z�U�a#zf�w��^�� ��<`�5Ĳ�bhH����S�gz�#��3@�G�2*u_�b���Tʦ�����qү۠�"��n;{����q��)�}B��֚�{ӿ��6��t��U]���{))���"�4��4�sҙ"�R��j�(�.*�!ˌ�i�Q/�1R��3A/Z����iŇ��'��9)��=)�{U!�ҝ��ڙ��~q�2Y<����_C~ȠK�Nq�^��|��F��G�?c10�f��o�?�\8�����G�1Ƕ�1��U�cY-P�_;s��?$>$B-�M*�k�lv���L�g��Fr2�s��^}\vG������0�׭=�P1�SfCڣ�PjF�51c�ʡ����T{�0zS�ό�=�n�7����y����� l��78�E�C�px���1�#ғi��*��4gGZ�0��@���T����2������s֑��r����WB���Q�%�qYJ-�$g��ؚ���w��(���v��
����/�"�[��<c��c����4C#;eOc^�����88��^qo	��@�'C��ٯ~*^�����7N�On� ��m]i2I�j��G1��z��$Z�t5��Q��ןx��m��1���Ęl�G��.��5�0Z��os
�)��i�sC`��E�f�j���q�ڼ~�H�Rq^����Y��.8��hκ+��>LTV�Ksv��@�-Z7V��c5���e��:t5����>?���'����"Ԥ
03^٬LO+���^#�Hd��<V���[�ݩ�s����z���ԍ��e�QR��עΫ5�Xg��?n@=k����{P�,�;���$3��}+S�s��wd�:i��$�V�l��e9"�ܩlK�u[\��ù��]�RC^����& ��Û��[��Ԓ`(�	<�X��sK���
Hc�$q]�!��C���h�JwI�^��_.1�$T�H���ǜ�4�6%a!Q��cԊ�k�[�J9��b�LW���!�׫��o��8>��k�oZ��z�����6�e�#ڄV��#浌e+��V<��N�,d�R�	V��Ґ��<`�V�q�'ޑ~\��:���R�&��=)���թ�"����;�A���z��EU�SV����VK��|�j�x ^(���ƿ/�3[4� �)�S�S�4Ӗ� q�ry�Ǖ b�sҤ��ێ�Aԕ���b����u,�K�g��U����s^��;��hZ���X���\Ly�v���ҫ���{b�������D���h���Zg��Z�>0��w��ws��%�v%Ԇ��9�T2f��*�����JZf�kHGjq�9��#���S9\t�sNe<��6�y�f� ��,)Y��j����b͐��1�Hr[җ�ڊ��>)�y�j+��$k� z�1�r9��z�dԲF29�0�q��L@�� ~�_h�t��ǁ�N��"��?΅S��I�������y�D�Б�S�����|��t�#P����!��M����o ��H��>��DR{ҕ1ƭ݌��UpG5�鹰+AѮ� 1Vb�TBJ���t��ܪ(�JZM���3=�?^��ܨ#x蹮sI���$����g���/���--�W+ۥg,9Q�a�x�%f���f�� ��7}�:U�C�*��v}X�)�x-���\��{X:�dn_x�$R����Z�����H����G�bC�f���S���~4��+�����A���;Qq0R $���D��$��68�k���`�� ��h��J���kȩ��Y�|<��R;���Rt���/���s�D>3��(4��^��I�N1\έ�:B���Y�#Ojo��23��3�9�"�O>�9�X[_��ާ[X�RH�c �\��FxA���� 
|��m����#cߟJ�r懶��2Ez-������H�\>���%Q+�� w��H�Ȣݹ�����y.���f�ߌ-�8#}d�m���6�7}��$ 1�\֧o�3�x��TM���[ōz�7�Z�Y�18�IJ�[�gr��m��b�ksE��_�I8�=OqW�C�[��{`���?�5^1ڨ/���p�#������տ�����-G�h�c�S�<d��!�5��xr6��C�<Wp��G9����w�r����$�b���Y��M\���sT�e�n*�6�%�-�꧎�՘���c�ܹn�4P^��
g4��};��Z�:;p�S�ۂ+�09%2-�y�P��NWm&�ִ屏0͟7Zc.*m�����N����u8�6�Z\mQHݨ@&�ڍ�s�*��Ғ����10V�� /Nj
z���4;�T�G�D;T��Zb	I�9?LR��Q;�
X~�!X�8⟻��Q�֚$�n��Ua����kq�ܥݪ1e9ܵΫm��xc]���d�Ғ�Vf����}'�s㐵�[k�(ȸ�Q^},Pź����K��{Q�ny����UF;�3|C����b3t�C�,��e��Ƙ�����eݻi$w<�
4�=i9�I�"`y�G��SH����V,�h�t<���mH>�=>^�R(瑚v�y�L�nOZ1��Jz�3��"�Rm�2;��0+/�;։q0I�ګ�Q�Q�9kK�9W>�叞����p��=^��0�@��7M&W�J��w5�ilrju�����6�@��Y��W����\H!\�N����cu�4�������_�� �Z0�z��P�}Ԑ`��ߥv�P��a,0F1�I>�x���g$&8����t��7^kQ֍Ҕ\�s^�� 
��&K��;8"�x�DȂ}�y*Z@p����2�ܜ��e*�j9��3h^F}�Dry(�q�Ԗ���y�WCN�^��DQ�n��k��o-�TIw�G5��X}�3�����xWN�"�]�95�ܥ�`�2�p:zW�jZ�ۥg�mz$��;I/������-�ĳB�(�H�s^r��Ҡ�s #8J��S#Q��d�:�Cv�s�Ҵt�u��K��j�^Ԑ�m��4�do����=<�k�(�p�z܍!����kMa&`�C���[}N�!�]��cU�B#��ڤ푚�4�6s^���א�8�K�V6Q�����P�ٺ�9��,E\��+dӭ��z�wlsN4�R%.�k���k���u�A�@�Wo ��X���{��Ѵj��c�t���)3��KS�&�B��jƱi?1�� t$�W�� cF�$�"��p8<zV��-6��QW(� �Z�]���4�lr�ܹ�'V�O���]�� �k?-TQ\=�up̧#5�`��.�o/j�OZU���/ˌ�J�q�b�T��*��a���O�0����Q�������>rx�m�җ�v7t5����l�jU]�ha��(��Y{Sv�zT��4�z�E��BcۏJOj���F�-�0R�(�R�K�����ӊi� <ӓ�b��P���NA��~�	|�4��M���R����c���S��ނ<��U&�TN{R��X(�l_G�W�84�t���y�C,�8�5v-"G99��CcEF[�� ���Nq�E*�{��4VX�sUFB]h��v��c^h�G����]|����U���s��G��8�u=��Gd���P�	x����,�eEs��g)�3^��ۜ�(�L�W���Z��(V�D���w�8�v e=;R4�LSy�f�q�3N=qF��4�y��H.0{R/ �F�p*�������������*��Sa��Fx�W�kD���q����Q���iw
v3V��.�¤X��3֛$�qڬZ����y�QU3HB��֚���G>�kF��D���N�)���~_;�in5 u�L�P���]̅ی`��=�1Nn�l�4�`e�x-����zT�v�Z�<Z��݈�5�c*
��RK�r��"�.��H���� x�+д�
x���_����>�I��݋��W��H����RC�q��z�2�F��Q�X�=~bEyU����&�������ڦ�������V��!�ߌ�;T�wg�9,ۏZc/�Y���"��DWߞԜF�
��H���������N��Z=��_Ĭ27sYX����6�x@���=+y�����O�5��Ŧ�����W%w�D��G��h�&�Ɨ}xY��J5Y����`W]���o.R"x'�ַ����Ie"�4^��������ǥ\��Xga#5c���ۛs_b!V�K.�I=*y���k���qz��M_Dj�����?qxC����Wi��+��'榿�]�T`�̿��V .9�Q%�GW�enD�ϡ�oZ�e��,͹Mkh~'3�#a�lw��z15��01޵K����<U
ԥN�T��da��NU����5��*�޷�3�ϪL$�V'���oK�#���j�ȋ9lz���5�ԗ� ��XS���V�BL��X�����$1I��N0+�4���6a����c�����n,�<A�n���;���/,�� �zW�x��Z�S��gA^Qqpn�C��E4s�L�o͚p�p��ۏz����4�qҀ~P�m�Fm��w�Qތc�Z_OJ��(�\��Hu�қ����QHx4����:�i��)m�}������q֠��^��G_��.9�w��1@\�4��{t�������HjM� �!P7zՅ��"�cp dgң�n.����㫱N���`�9�J��4"��2MY�߇.5	��"Gһ?�I����xX�����B����i�\T�J��V�XH�\�-�c^k��w*zhSLF�c4U߳��Q���*���*GZ�����^��x<+�A��l�f]�vʢ��8��؃�8��GM8�z���ZL�U�� 1�c���tӓ�0���*�l2��z��Ȼ�LVό�7ӯ8S�ȷo�����xuW+ e��7b�h��{Z��3R#�Z���K��>�2��ir�0���b���j�i��#�;UX��JŔb��q�)�g�-Y7֜�sH�I �Nh�:���A�ߠ��=�c9���6&�m�D �ԕ�i�5�-���֥�E�y<Sn.1�͞c;arkK��E�݅Ħᶩ�Y��ڹni��������BWܩ�˖ ��1Z�6z�r�y�k5��0Ha}Â*�b}my����1��.��5�� 	�O���W���fp7Z��^3�+<���c^�k��j��� ,�5��Bzu�� �z͵蹼"�8�ؤ����H�4�"<�R>տ$�%�ʤC�q��^a������12�:��-�s���ˇoRM1�q�OE<�)L�7�$Z�����h�c��۸�b�q�]�{�m��ٶ�z�_�&���v�[�V��%��^V��b\H���j��֬���⽽K���)�����������
��3R{�RqOԵ�."�n��>R�ԙ�u�5�s�gK!9��J$���T����X�覈X��Z~�E�)c�����sMI)T�A�w7��uog`w�#�9�5���������XuqB�g�������q�0�Etr�S������T"�|aOz��V���1�����{�Vl�Nư��.�ł�+c��ZI�WfK(f�<���j9q��Ȫ��dj�R4���+��}�5��%����{��$�s^��];Qԛ����M'��m��t}7M�H2�ီ+����y7�������/�o�����N��7'&K�y���1���	�4�V��r��^}`�|̨��=kٵ�Mf���c��MwI��.g;����FS�2�d�R*�]���yg���s�'Zw~� 9�v�T@c4���1��.�1�T@m�J���QK�Ոn��4����������K�Sv�⤻��4�?)��<�;�\��J�q��)ξ����t�!=9���ri�~n*X�=��ђ��1ޢ�t�5�ra��Ԍ� �'�w_t5�|P%�d/�rb%�ua��#޼�;}>,ƹ#�۾�V��	�W��v)mf�v��n�.�����F6G�z��6�F��=���<���)#>��n���"s\N��T�\𬙴]��_H�5#W�j�6��)h#�mϐeϨ�n<�-�ʽ*=&>Z|�Z�g+�Hѳ�"�ㅰc��i��V�qǥtچ���N�sU.#ڹ��3]��ύ"�p?�y]�PZ���fb���^I�M}X�.)ٌx��Tx���s�G�^���m�i�x�m+�=��;qO��(�)Ư�NQ��A�i$e�x�@�bI5JF2>4;4́V�mNy�S�6�
�u���A=jĒԚ%�B�&�����Wu]Gq.��UF�V,�v�ph��ۆ'���ہ�8����Er�>�N��#�I�dv��mhs������ l�Hs�͊ehxu�=Z~��\Of����4K�D�Ld�
���5���nn8��b��;G�!?3G��+���
�˩M�:�Q��#$Vz\�m���N������ūG"�7���|�)��H����*+���r����?���HN�L�>i5�h�����*n�J�\��1Un���>�����V�����^GL#oy��ۙܓǥh-��MKZ�� "��J)nL�s;""5�̼����S]Ϲ�Q`wr>j�GM(Y]�l��sC)����rz
�O<�+��ٶ�_��5���?�Wѫ���ɪ�ۙ9�t^c�A�l`�x��>�S�mC�84}<yh��:�\��6X�+p+�}>KK�Y�v�^;�i'O��3���099���A�b_O��ϿJ������m@�qҸ �jm[X���\*rźW�x�춺y�'Q�w⥫��P�wR'�cClYw�w0����$���Gdd�=hQԹT��+�%q���χ���Z0�d�^Ou0E�#9�U�sun���ltjݖ�Q�Օ|M�
M.��c�Ň�=Ӝ�I⏃����مE>��d���~ ��	'�!�B,T�Ǘ��~�1���)-���]�������x&��ǆ2�&�e��>����a�/�.�&R��>[��4��2�*�_����b:��R/L�uFɥ]I�U��ر�sI����(ԞjD?�>���}��X�͉q�4���n�ZAzh���*�9��U���עi���UZBr�ة��=�R��J��z�8�g&�O�D�S�P��zO�n���lx��_�Ľh���S�f����K����kEla�(�
6:-!{J}��}&})��ۓZ`CNk4U#�����c �6��a�fnI�k��ރk|�z�Ծ$�7ٕ��\�gh��5�$�9�p͚��{�m��96��ӌ+��{���\Y#�Xר~��G��	� Xr?J�B�d$c�J��GL�Dj�Tv���lva_�}�Ǻ�v�qO���`�	�MCO���5�uj�%M|�������0��EQ��Y�����������(���!s�����yT�ɬQW!j���i ʶ�j��#��Q�j���o_&�b�N0?�z.�2[ۼ�6�J���׎I<J�>p�֑WvFS���� �u�5F �}+�Q�<qڮ_L��/+���U���{�|49`|�&|�+7���h�a���e�a�sK��1A���1�E �H�D�W=�@y��5�5Fi���Y��v��j�Fk=do�5v2�� g��\�Qn�қ$��Vu�����qޞ�!E�wcnfi��mf�)n\RZ������/��ݎs�刭�^���P�M%js�}qH�\�Q@���9���H�(���l�+6�Q���V�`4���O�_:�s18ݽ�f����3������shߡ�b�J�f�¯�N1���oG�[�U��P�^U�麅��P��ā������[�]%V�-�&y��$�a$��I&<�W�x��\n�A��Z���B� �5N�<�c�I��F6\�lV�#ÃZ�±���{����֚IΣ��d���I�ڳ.�����ww�#�j�U��jtҧev#u���i=�?h��)���r:V{�C<�����Z+|�f��v��V��8�M@�um�"�\�N�1�a֗�	�+NUc��:oL��V�cޱ5+�r�^޵��U�̍Qʣ��o-}ĭ���̞��n�ė�e�#�k|�H⭪�9Q�B��.RQ����*9�X�$79�Mr���޳�L�q�M&�&oV1��]O�f��d��6���}ku�0z�+��N��p�9,z���h�G�h�����dsk"�Uɫ���;r�<�m9����K��3o-�=���6�i-� !����P���P��ޒ3�n=1^qto�gw$��{֥��/[5�.�62�+üe�}C�:��wY�����Vђ��.TwPq�b�M>^Mc��r���'�U�b=����#�ǵd��b�%R:�l�rA��/b��tg?0�bvj�����n(�b�3cr�jU��G�k!Zv���#,ۺc����خ���B�'�#V�Yg�A�"�&2sҫ���ǹ�n�f�⏴/�d�2�ʮsH�N�1���=�{�� hNy�-�|�ȒW �=i���}}is1{�5���'���	����e�Y��o/a���f/c涛�Ig2�M�s^����v�N���WYl�)*��ֵ4�M�d���Hvp���W��o��y���[9�6?�;G�#ԡX���ax����Z.��q����I���Hq�U���P�x��I�Z�5����`pEu�\q�/m��"��DoNG֟�!Gqe& rk�-d��=�s�W��u+��$��TS��G����&�8ndU~��_?Z�L��TRG�IȄm�.���ⴴ�iڭ�:O�#p�f0Ȥ�\b����\BW�t���&�u�}h����ZNӋ��+���s�X�\M�������{��{�s\��PԲ�F%���7��h�=��oƅ���ñ�(��z��l�f���C��/p�܅��n�֯k�$����Hw���V��ݞ}\F�G'�hmr��oC\�;�&�__Ip��z��[�׳dy��mS��Z�\f�]�4���$��q�P=^�3�-ǵg\\��(���z��ϝ���vGLb����KP-���RH#^}8�f.H�nn7�N�����Ě��p95-���
,�y�=j�6��q�V9�G�A��qLf'����~���2�(����6�0�y�s�4Rc9(�� �-6�o�n\��z�׼=�J���6�k�xo�-�*9��d�%�2�u���k}U���E
�m
��(�T���Ɨ!B����򽟋��.�q+��'�85������X���Xr��gF�]�]�۴ڴ��o=jXm�X=sɫW�&��Aј����2�:����<�sh�f�Вy�7FE�ze��y�ۺ�I�r5�%��0'��A�����Q���:�8'�*ͽ�q�[[f|1�Z�[�#��Kh�c�q�7��wZUQZcy�n����=��*�x�qw��ǥK4�y�ۋ�́M�٤l����$3z���8��J��iO�Y�6�t����������I�6azE�F�Z�ko��8�O��������ԛZ!���Q�s^H!�Y��Q���
�𞲚m����E)y8;]�>�?����ZI�0���{_�+�wU
>�QH�$��rOĵ�v��`s�
ܛ㴉k�$PH�+[��eƭ�4?��۝���8�֯���{Տx�}cv�ǚ�21f�[F��)���.ޜS�̊�u��q֎sַ�F<ϸ�!
�G���T��9P���/�1�u��G4�Ps0ڣ�
]���S�H\�s*v\S<��Jz�S�K"���?:,�v	��2E^H�7 ��VN)Yt.�8�XUI�U��ަ\m��UXs]_�.�1!~��r�� S�����y5p��gu�oë[�@�����}&��8�8ֽ@�"��f��rj_h0�6���ʑֱ�ܤ�8�?R{Y����z��èB�-�W�][ͥ�c�3��]/R{VVF�*���Zl�Y�4�-<*�����e���#i����owg�pq�+������6-�KC��R��9����N��#�3>���O�e��*�W����i�+\��t�z��$iJ��+��_���w<֮����5�}�N� Gb���?����MG��z?�G3�Q^����[
Nv��1�OC�G�^|^��e���4W�ū4�.�)}M<Sev t����ϕ���e�|̛OJ_3�<׶���r�SA��0B��>I�f%�I�4�@�Ě�+!]�z�0�y8�C|�b���bڞ�6i?���Mf��il=�;�'�fMp�m�k���j�ڬi�c��f�Ψ�A]�-���Ú��!@>�5�aSڳ�.ZW;NI��Fvu�����{�[�E��9��5yT.GC�hI��.U�Wj�8��ך
�\g�ס͸nE��Z:�Z}ăzTrةm`�8�短B�nƎ	F�$�i)�9�"��tj����@�iv��@�G=�j��xF�x$�NY�s��YSv7�E�2=�F8�˶�\Y���o���U6��Z�\��2N2�"�o%	�k6I�v�ڬ_\	3��}sL�P�d��e'�����!��v���kF4ؠ�C-��*�MK�"��N6F5���cROZͺ�,H�ۂ��N�E���S���*}X��B���/=��:��ڦ����RCj[� ��4�j����jO�Y	ظ�>�~��J�-� �i�q�J�ԓ�Z�yy��Aމ4��'����h8��� /@п�#?ZKkS3n@���f����)(+!U0��t�HaRx�?npj�Ld���\揼ȿ�6p���q Ebq^��~�7?�珞�{�i�ۏ�HN2:~�U�w�O�$ǆ�?M�xSZ��.�s�s����g�啙�C
��~d��<?6Cg���i�eU9Bx�y��m� d�_K/�*J��]�q�3��}3�p�
�,[�'���b�X��g,����ْo�J����a����W�^����m�Gߖ�����Z���� �_�3-Ŵ��f,9o��+_W�l|gq�q��8�>_S��3��_Km�v�+�pj��kզ����p���~ju SJks9���h��m1IK�(��Ҋ( �'�4�zg�J��ԁ�g���~�G5�l����@�dp���_z|	���)�xvդ���G�3�"+e�篽y���9X��QN	��(�������7�=M}�����tˇ�O�������+�_ن�[+f�z��?\�\�u�V,�顐rCc�6�����,n��C_r�� �-��C�c�G`�B��N ���� ���Q7�6������3���^w���H�b�Հ#뚻Z�/���^����3[�|��	����/�V�G5��b�F�����^���r�.֧Ƭ�OJ�q8c7��|?�lY �=k��m��nZ)T��:�{��sqX�#�kG�5��c��&8j���R�h��9'�u��YX�"��[�x�	��1�QY��p8��3��þ1�{��E�H�8�&�g�+��*�᭄�}��}�����vG'=놮!�v:�ᔕ�ę�7yj��6U�5],�\G�}�����<Os��#��Oj��7�.�x��p�g��rc��tKg����)�����?AS��������.fgr�H����o�)x7úލg�[-��34�$��X 8���z��m{�����tm7M�m��������9?��<S�?��F~E�w���"�:��]�l��5����ݾF�2&��8��S�Tedy�ͼ�77�8����&�t�l�<b���
1]����j����(��'"��5���zҳ*>)�A�4;x��:�F.����YW
L�>�7�kܳij>��j��~��|�j�� �����b����ɩm,^?�E��Ty��kB�RX���y����b4�Q����e�������l�z��^��_��:՘��d�ݷvi̒2Qw��iz�rL�Z�4��� ݟ�l�C���2�o-��S������x<���OZa���c��N�y��;���U?�I��_Rf_M�S�Dr#�ZL�
#�q�E{U���
lb��O?�[����Ж�ar����r��V�^#S	]�A��{'�I3�L���ޏ&�[�q�����ݛ�R��<��PY���c�_F��x�5�p�Џ�-�>O�Rx����yfrǶ_�w�VA���|�&m��>��cg��������B#��N+������°���#�WvqB
�����|�r�Z�y�C�֩K�0�A5NY�F9��S�z�+n�zSF3J0��^��c�<�;�HI��V-�����L������q�T��I��$�1�Sڒ��y�؞�.��q��{�pX�*�������a�L��� �U{[r�'�Fe9a���#1P�6�J�+�}��r�cڒ>����z�;�5Է��K$�S#��i#�����|Yv�X��|py� "�K�O��:��%���Y�n�l��_�3�=���;� �}��4��G��]�^����/�ϫ�RI������V9�H��A����DE����ͩ[xl��l��^���/Ƕ��n
���:4k��_���;Ss4��3���W��7�أ��q*��
 ;u�A�'�U�f���z?i/M�5�n,9�kN>�'���Z�7��Ę�257����Hv�橗,���~|�+���6�\����9D����P�ގ����� QE
�5<Tt��i���w1��[�nk��g�Ě~���z��Nk�9_��Ǯx���_�ȁNJ��o�s�p�8$��Y<[���� �-����8�3^S��}���溭�I4��q�yM�z).���~��K���h��n����V� �o��J����
ɰ�u��ZC�Z�_<u�z�?�ZS����qN,�ާ�?�W�f񯋮�f;�1�ӓ�y�ɑ�*�i���-A9'� �^o-���m �L
�L+�O0��5�H�4�RW�D�W ������+�3�޵�V���F��
�Oʧ_ZMh8��c*`�]V*�������~#j�Ž��=ԏ*���������Ǡ&�����W���>�1��`r��q۟S��%��ȿ��?���SE�[FɴpH��\6��?J��J�����W?7�u�v�=),o.��v��a���#��j���4�e���Du�(pE|k�{S���9����p�95�G�����fˑ�W�~"�k�yUy��ԛQ�6��������Dgh�;s�ڊ�����p�;y���9�O�~;iQ��,��mٯ,�~Z�o�׆k��Ó���(�5�t>|�'�$ ��LG�Y����a?y�u�����R5?�5�t�h��{Ԋݍv���(�$����.��m:ᡸB�8��̮#O�Y�9�z֥�_J�¥�5��|=Ԭ,Mۮ@��hڒ2-�uSP^�55�YJ�4�7(�n����'�GI����N=kI��_�* �]������я�$��|�t[S4r��%�`P�kַG#������·q���=zm'@gI2U �9WϺ[M�\�ߎ}zW�5��e��b���5��;3��<A�O���x{K�Ԥ���,=�]�����Ci���l�cdr�Ry�~+�?c�>O�����{�$��'�־��խxk�z-,h5W�ۑ^\����=,|/o��ű��q{mj>��� J���Z��pѼ�9��Rݢ"�#�W�e��|��Z���To�� 3B�\�a�9�i�G'�j�'��9��F����Bʭg!��?�V�G�#;~�!l����#�"�:Ưq�F$���R\kڭ�ލ��u����������}�� �Pj�8�hVBW'���YKgcx�������ƥu��~�OJ��񏊴���y%����#�NA�������-�(�G�K�.�q��5�['��^����:�Up�6��	>�~����T��
��m������[϶��vU𬏉���<��e�ϵu?|Ea�O���[�
��@�r� ���*.�z�2���dxB�O���=���M���=;o�y����:~U%�&F�jXm�7���ƪ@"�#�-��=�7�R7�F=�W=�V�}D^���y<R1	�t�T/.����R�*1rawt� qP�۴�#��%�����jƢ8��P��ΉISVB�
ƀw���I��s�]�kc����]��=E*�TK�p��F*e����=Ӆ��t�-��Ď���<UJ�@ܳq��𷉴=;��Ɗ�8^���_��7������t�_tx?A��E�y�?�|~.��K_NPM� ���KPͳ�@wEX�v��;!�mҞ«�v/c~�s�Q��3	<��=��+��K��u�M�i���ny<��Wㆰ�$�Oʣ�k�/<I5���ǽ|��gZ��`�9�EuQ�4�0��s�o&/zǱ5:1��:l4���#/�}�����1�w��LQKǥt��Rb��C
(��Z`%I��Q��b����������]� �y����@��#�{�G�u�p�&�a�_�X�5�枩rG V$��>ĳ2��
���j���	�鮠�]�s����Wf{��qL��/�:]J�-�nk�������7��E{�B��>��v���^���-����K�bY�!b���x���1�'�s埉
u��Mqs5��Ē��"�sWQ�����G��=�r0�+�٧3�-�_C�Uu�y9�RZ��f�v�\�>��� ���[.�{ՅmVU�Q)#��%�LV�ܒ{W�|%�V�|��Ac$�/?(�y�=b �C������ya��vW��r1_�V�2>�jh�]zk[�m.�e 2����7po4�7�U�%��t��'�9dΡ�))���q�o�5K�8�/�%�����W=ob��w�.5?k�V�M��9��G��״��ĩ�m�����íCH����Bh%��K5|��ţ��<N���?<��a�e�+������c�M�U?��0pAZ+ю��>���� �_��W�G��
���V\I5�Ȼc���P�����<	�S8�W������� p�~��J�75� �f����;da�GM�A�����,LA=6��ߊ>�R��l����*߄>
�<�uv˅9��L���.��5�q'C�Q�dS��"�U�(�9��Zg�8�B���ڧ��%��͏lW�x/�X�q�?%���Y��%׆���23�J��r���y3Jf5�i~6�D��^��:\-���n������PQ� n[ֶӔ��S���W��*�ߨlW����7Dt��B��+#K���V��9 ������w������+8ŶT�[���ě�^<��ӭ{����!�
���W��L�Fگn�����Φ���&���]ⳤ�HQ�͒˟�]G�<m.��?3!��x��<+�:��+˰o#�J�/5�K��dQ_;Y{ǽKmOe𥨒�� �c�k��)I��!#y��D�_��L�]`d08�&���Z�j��!{�k�;�hZ���n��lO�����-ƕ<R+�w��� #�N��I�Ɗ�D�p}jK��:2$��=Aѡ��u���-�IC�����_R�>ck�'6~9������X���ᙐ���+�?���xh��f����#m,r:���t�`$���O�j�^��.�+���=+�|Q��J���~l��ܽ��Ѥ1���n>cUܚ�G��u���K�9�9��ⅉ��.��ֹ=R�.>I��U��_�Gd�p���y5-�x:�R�ON2?
�L�1��b2I��(a�Wֺ�9�NáO/�S�nc�� Z�4��j������,�Z2�pEP���5-��&%����V��'��RA��V� .J��:%%MY�(f#ޓ�h����q�9W�Eڜw�2lJ�g�NQQ�sS�y�j�@���̄�EJ�wqM��"@'ڦ[O�E��GOգa� ���<x��".�6�Z���v�훥M�<W�xz�[;Uh�+�����k��>��m3R	<���
˾�4�>����^}�˫U��mޢ�Z��{����O�9�?�V�أ�L�/���P��^�;OkS&z�k�<+Kb0�ݎInk��1i���y<��z���h|��|��x���'�5Zo��<��X��}���,E�����F+R��ns����M��	E)�% ��Z6� LT���{�x�zr�im��'�^���R�˼F��~5�M�x�kw���^���]¼,S>�
��a����yW�h7��8�Gּ_�z���>�G��֭/��ܥ����Y�����"�Y.��\U�%�{ذ��zF�k�̸9��y��"�ޠ$d�+5�g�|d�m������P��ǿ5�?�+��zt��VX��|����ϔ�:(���{SLt������1V�[���qҨ�Vmr[���j����
�Qq��}q�4���%�e|r:��T�i5(cP���5�7�� �w]�쭮�ű�dy����_�Y�}�_us��<e���wvO�W�����{�TG#/_Z�4��V�Q!��֫j�	���یQ_,�c�G����.ة�S��ם|n����5a�2s��?�}G�Ꮣuw,�ٻ,@�+���cM���Dmoq�e�}�<�S��b��;?���D��ʊ��e�G&���E}v<��>'����ߍylw��& ���^Q�����|�+�:� ƿ��X(��>��מ2���,s#�I��-���r�6��:֞��{�����cNp�fp������տ��Sy�x���K���_6���\��O�ɹ\���kj0����wg^����O���U.�=���jK������.�]�xv[o4,�1�=+����'����5�/�40���i����sJmW�O�:���[�V�������������Gۓ^u⿉�,������ŗ6jU��T�q%�[#����).�I,���ݎ:W3T7%�(��P����v6����"WT�O��J²���sA�\j0;�׹����ۈP��_�
�Q��w�������� �׻|6�Y,�+�IF��q�Ts�niʠ�>i���Я�#G�3p*U��"�7;}+�M{ᎅ3<���6B�TW�?�����@��Z�-Yܫ�O�|M{K?-�G�3�^8�P�%Af�8����Qὧn�'�����>���x_�1Y}]t)W]O�!��+�I������1��{������M(�� t����E�#�#�R)}\XG��~8��v�׵wv?.��1.Tc����T�%�d�jG�v�� �Z�q0� �
�<e3�)}\YGκ��澼bL�S����Z�e��k�X���"�#s��E�I��I�o�f� �[F��.��>q�{>���.	d��Q�^��O��2��U~�u5����� ��C��n�W��⶙��4vZT�;��]pz�U%ws���lONr*��խWAԴ9���4�8�n�+������J2 �J�^�=���\*��K�q���K��
��V��9��N���a�ƴ�j�Tnt�J���HW�f��c�9��F[5�����;�i�)3I��.;�ɡ�eF�m�U�'�Oj�$������?
����N3Qi�f'�������k�U�Ψ�V"�a��q.����Y�_Lf�F���&��W(�F�R��+q�\ q�׳i�*�Q�������ȥ��;N�%�V�H�	�ؤ�#�(�i_��.@�� \q�s��oZ��x��J���Vq�q���ٳ�����Ob�n+�Z�>#x�K�d �d�}�Ő�ڸOk�^�1�ɯO
�78kٳ�nn�\�ޤ�sm��/�1�z�i���W�S�����R��?ncߊa�5_�o|Q�v^�����{"��=���?�A�RI��B�H9�G���]�#P�4��^Uk}��<S��g��=�����K���f���q��Bm�A���f�q�~�=��Xk�91�Gx\���e"��|1���\^�v'���� ��&��'�1T�����K�{����^����r��(ǕX�]M��E�nfb�� �v��+FiYV<�p�7�[8����u���╕�򓞤��+FNZ�6�v���s� p+��.&����|�sK�|L��\�Q��s_�Y�ė
9��J�����V�6��� ^��|�[�i�{�� ��m*���˛�#1Q�5����<�RSV3����횑dUdc�����Sv3^��4x�rC0猚����!݌����p&�wr0j]v��qè�by/L:���wm�{f���O�P���C��
���W�����<��W�|6�垇p��v�����/Q�A�J*����^!��8(�Ҩ]|J�
�����kß�١TP��^k����}�;��$9^k�����M�|b�h�UϘ��W��L�ީ�fg��� 6{�״�:������-7D�����Ӛ�����Ril��L�#�5�B�=/�M��lk+a�����E֮,a
�@�W�
�El�6�x��L����N?*���k�~<F#���+��z���߸����B�T��zҏ�G�]'�Kri[ӽ�'4��."����f^g��Z�n�o>V��Y�cz-ܳ`7&I�_g�y����L�랕=
�c,��֕�ۭ�k��8��Y�4�==�J�=��#��Ml�ϡ�-�����,�.N��Iw��L��%�Wc|��+3AY!�Y���׋cO�_5�-�I6pz�pqJ\�u*~������fу�2?��[���y	{���x���~� �3t�x~�U�5���&�B��C�� ���|;��ͭ�$���p3\��E�3Y����|uI#F��'����3YW���[h�ݜ���}+�<Yb��N��d�1���m!�H1 ��5��Lh�n{%�ǈ�����0*���v�Ddz�͗$32�d��K����jp}L�sh}'��#v*UF0x?M� ��3vU�� g޼GQu���_1:�' �e�Y髤��vӪ�#�?�g���b�=*O�ү.P��㊫k���9�>`��s^g��}:�NWp�+����y����(�Ec�a���4�^1*8{��.?���YK0�1Z��к�ϕ+!$d�9=����;~�>���_�~]��+�d@A�޿3a��xg�7�pQ�L�ⴥQT��M����p�L�F�$��3^0�Oֽ��ȍ��~�`d���.nB��^s]�zn.Lm��U��Um���na��ғ�y��Ԇ=���(�յMY
�}Fn)�2�'�x�ri�in�!�:��I=X	�����j$ri�)]f��key�j��q�TJVFшH�����\Jx�R�'�q�=j�����wS��hJ]TGsSj�ݏ� UR��h�h��ѬLK(^��㩱����������k O��N)	\��T� ����.�yU˱�*H�5v?N�88�3X��p{1O
�QY��j��f�x�n���jV�4��[���n��i���銞D>ft	�y�;q�T7:��|�񞵊p�P;Rz�V���/4�?��TM(�Pd�=*)��Pj�ɲ/�1��	3����K!�9�~q�sG3�.R�n6�F}�o<(��f�R0OL�yŗ�99��9WR� ���c>�Ɠy�~5U[����Y\v��Õ������v�Cz�!!�p})<�L������ʋ�i,��_Zi�7=Nj�����R���>f�-,�y$t�%��j��Ó�H� T97�I#Z�Z�6_����֮��{���V*H�0H� w���y
�f�q5�hԸ��/�n����y&���
�\c�*O:>T���3jȻ����P4̼0i��>u�ߺ �"���b7܍�m�=�?�q���4j�,���ǯ�W3'��Ϙ�b����ޫC�d4��7`��.���`sNmFK~U����k)d%�z��e�r��jj����o�>�<Ak�q�c��z��<�kg�ۚ���ߎ"����b�⾕��}v��E�򕹹���k�,��b���0W5N������
�?��#m�xf�"�_����|�H� 8�U�ƻ�?�K�xS���� a��|����=HWPn��c!��_�/�F<�X@��_�a�|+Il/Z��^p?J�a�ɫ^%�@��"�wÿ�.�&��Iܳ�[�$sF7W<Qf�����+�[OxOR��[���`��>���76f&?w�*T��p8 �G=+*�1�\�Wa�� ����0���+]ߊ��iZ�*a�L� ��JKb�Ǖ���x晩>ъu���u� ��?�[�j�n�V�͊].8�|�l��'����`Rv�½���]������êg>�㖶����"��^��hr��{�����m l BA�+Ǽ|m�t���q�S��[K�oȸ�ǀ=2+��c��� �\I5���g���+�������+>��o�F�vդf�'~��ڳ|n����e��p���^0ccj��(�s�¤�&�5��������&�CԄU�Ϋ_����!Y~��w�����y�>�hSJ�Jp��8���n��iraHC���yo��G�Fpݽ�R���isT|+i�ܡ�rh� �N�v6���>g�M2�9=3\ʴ��^�=�I��ut]��x5����됈���:��&�o^�	�3�ҽ���"{,����L¬R3|U�4���}:�l�`�w����V��Gڙ�s������ ��;w'8���Mq�֥�OV��]�sJܶ?@�{�T���y���N� ���5Dּy$�,Y���oy�{]���J�t�A�(���5�a�J�UtGW��]	��'ڼ"Zi	�_@x�x~N2>���l��ҽ��{�*b
�)�����Kpkmˬ�v�ȧ��rsP��w(��l|��B��rsȤy:�i>R8������\+g�����zRɻi j��̻}+�R:�d=ON�ZBx�&��m\�uYɐs\r����:D����P����O^M/��B�G_SF�Ť�����7*���gӵJ>��E������J��|�jg;�(�`g�9I�������Ӑ1�'4�~n�d�h �n�.����#�jh�-!r� ?Z�M���>�pNj��Y��|P1���9�B���#R�u�4�|@��S�>��=P;�>D�4�����F=�NRJd�Z0G\ӆ�2x��U;����2w� ��M�W<`��3{n��|�2�=*&Ϙr*q���>H'�(1&ߖ��<��:�0y�T�Wr`pZ�����1�w�_�Z�ւ�wV��q]��?[x��Q}�n S_��9�;M$��4�yq��W,���#D�S��?��rl��9�M� ���<�oc_���_��9�X�)�Cï�(�a��O��SE����ZʮM����8�g�ιȂo~9�ӈ~�A�2I~���o���;aO�/m.���*��R�P��"��Z��i�P�c޾��àxf�9a��׀z`zW�ڥ�ZjR,-�g����I�s).ţ1S�H���VUe�nI�R���� �#�U��@�8�����R)����[]�q�k�l��Z5>c����� �u`�"�Ϧk�4�EŪ���
�W1�SzX۸ק�O���mF^���Qh���O�湬���� ۗ+����KQE�]�����}��O��A�{?Ǩ� ���>я�x�9�{���o��_��3�ݪ+���H��/��8L}���ᬂ=Pz�y�F��
;��$����V<wN�e嬄��}rj]C�S�jI�<��a���jy0F��������otxD���kT�>��񕽚���WU�]\j�� p���"�C��=B02y��_�2?�n���@��j��{�
�:�+�� :�/ ���C�(�(l���\���9�V�Ḅ�%��U/�Q�9�׈N��:)d�ʾa�ԯ�J��?�s�Do���u�u�w ���sYGC^�����	$�}?
��x�-�sa�7��k���e��HI���}�x=�4�&��ֹk|,ꢮ}�x�5+`7�w���(���W�y�Gn���z�!~d�c'��kĒ�z��ze�c�F� ��Q7���^��l����j�ui��s��R�:)�Nd0W8� �<�~`l�����k�=���rIϥz��.#�f9w�{Y�R�����r���w�q�vQ9+����2 �k�ZU�R�7?5{��/4����|��k�]A����5�S��M|K�n1Y��� ��?0t:n�&�.I9����^.�ӱ��ztJ�3��]&��~Z�fc�1��c�#��H�ˏ�׍1��s��։�KPf�������ޘ�����9��J̓Q�lTJ]��/^@�,�-�j3�XI��#[�Z�4�GZ��k���̘�Mqԗc�����B����ŵA��i�ۮ+8ǫ5o�:bP7�CI�(2e~�=*����U�]�����(nR+��JT/$�`)���=9�\��X���4����#h�зL��,���ӽ~�;u�c���jO,�B��hH�նn�qP$?*��Z�h9��d�p}�=�#��dn�
*�:���I���Y<O� ��^�׵ *�)Ȫ��¢]ʼ;T��<�h��_�"��ʚ��^)�B�=y�@�C�C`�U�}zS����
�J� �c;zf������zTe�|��4gw��U�5� Glp}�����w�6��1I�����Sx3WI� ��_Ni?������=k��;X��K���qL�3Kt}��@���g�j(�;�A3ξD]V�z9�Ǭ\ ��5�3_h�c��	p�?�cj_��M���_Z�`�Pɨ�"��	�٠����<��5�$
۲pNk�`�7R�s�{�Ab�NkOK��������s���VE$�6���e�Fіj��4�V��D���K&�B�ޙ�#�����V���������:���Ŗ9V�7W��V&8@� W��?P��1B�B���y��k��?y��%��	��/�ҧe=���N[�8�[��(�Wފ.9���$�<�b�Z�8�l�����pد���ֿH���<V�/i:��A����񥞣
�j#ͅ�k�e#}i��MjAG*{s[�)�񕏨R�V�[X�M�{ W�|E׬�n�eY�d�E�ð�@�5�3�ě�l��Q�[�zǀ��� ��H?{5�����ɢ,DF0z��J-N���\�1E׊�q�v>���)˘��xwñ��iȊX�+��d:U��أe�Fq\�kW�;��5Z��XU�sڝ�~����o����+���+Ŗ~��1E�n�{�k��?^}�!�Zvz��]Ĳ3$V\�M���icS�����|�yu�\9m�~�����U����,����2�O�� jO2�~s�+�����FI�B�j7�A]��B��<W�E��� ����U��/�����Q���Pgz��u��I#�U�kT�)�g'ּ�I��b�N����5���[��C\5h�huS��=0\(��)�jO�
��I�����R���U���
�����n�XK�Y>V�f�M\��2��k������+�^���=��u�N�9��L�x����1�Lו��������𮽨���Ǧ	���_����ƬNX�^�:.ǟ:�ԓ^���1�������b��@�[�u�u�����8���������b9�/ ؇�O5�N<�<����$��0�,?�x�l��{������T#6� ��3�7~y�NCȖ�:c{�~}�Q�g�ꄆ68�Jc��>�Ӟ��L���j�����$�>Ne\Hev��jKKt���dJ��)b�j���J�6�ӵr۫:�����Ҡ���N�n0*�V���S)v*+��x^ٮ$��t�� Q�A��j/����Nׁ�e�q�Z���(mܠ��(�#��5`�s����R��_j�ؓhE�j&`�<ӕ�0i0{b�ɓ�8M.���R:�
C�?��`&�_�H�����b�K�����2sNM��b�3d�)�\�fU�s��YT��>���}酶� ch�S�y(PZ��8?� ;p���u�.y�5A݌b��h���h�Q��֓�9�� �W�����6x�����A�`S�z���[� U�@�zSY@�@g����ޫ����P1Z�YPX�ZE��9��Fe� f'#54zJ�7�_u_�9�y��pi�.@�4L���)�����¬y��qǭK"��798�As2M658ަ
#* ��@�ۂ*<I�9nON��^��i�F)��Ҙo��{r)��@���<��r�V$���R�n�A�2呜��}5]mF}3^?��oh�8�m�*m��^#�g�Kav�y�~\w�R����{�z�%�ʳ7����*iaR:��Uq���
� ���R1�z潯�����1!�_�k�#��_�a�|+�G�I�riz��X��Qè��Ӊ:f���K���t5B� �Q��ˆ#��g_d�#����Y�[�RjM��yi���$�Qе�i�y�=}M]{�j���N*�����{V���eę�Q��/��</�J�M�#I
�+�4���į,�V��
[8a�2�'&���ڤ1�k��&e(�mv�i�k)C}�N
��UN��Q�`���%�5;��g�E%̲>8�Y���h��%^��WZ4�}���<08�+����ک��4��ͼ�A��N?,��C�v�FX܂��5���7״���c���\���i��,㏚��2�
RL�7��Ą�«Ÿ� ��?J˚���;�~�:�F
�����W�4����|+h�,��0�\WK��:l�V9���
�����^'�n[��l�Ғ�5Q�OQJRkC��a�b�@�^��en4�W� z�y���_��*ZH囧�v���>.��M;�'��I5��FJZ��6�4�8��bǏ�����ɡٵմ�︚���o�� ���]�� ��B��r� 6@5q�d�Ecõo]ꛢy�{�5������P��ޣa��J�{�N���c���� �3AϥI&;z�m��f�6L�|� �P��I�j��W�M.�h��ȏ��ɮ)k#Ў���cq2�� u�rHa�a�^�u����(�Ҽ�V�n/���J�ES���}�ێ�f%�S�sL���-��d�U��B�ݚ7������6��`U-8#�Oz�fwq�
�����j�NjL��S+��R�9���H�硧���?
{7V�J �"���I��x4	I�XqL.3K��j��n����Hy�zX�l�d�x�i<����,1�Tn��i�f~����Ͻ0$�� �z�OU���H���(2ڐX*�s���]�I�T�j/˜f�^���Cs�ҡ��8�-&ь�}h�0�x�Ot���`�Oz��� 9jM�q��v�x4�	6Nx���3' ��V��v*,/ i���˜б��Υ^'��w�h���=}i�e8-ךFb���E"�?Z ArE5��ޟ��8�ȣ�Ny���g�5s�R�z����j�x�sP�2��<S؂G��9�mf�I��G��?%!�={״i�4+�F+�|��x⽟GP��^��b7=�[� �Rs�J��N���Xc�k����ǹy�O3��EIG!�E9�K�W�Ǟ�~��dx�A��9�����+��?����|bH�W��V߇|��� ����3�\z��R�Oݯu���ֆe�B��#WD��a�]�c7��j8�$ѹ���xwP���;�Z>xlq^���\��yK <��S<u��?�^P�	���*#)_R���Q���i���3�ֻ���{]ygb��+��q�[p�7d;@n��>,60h/"?�z:Q91����?�fF����h7� �˴��nj�Yui�`⽛��0��!�9���ޅ(��9m7�-�B�Mt��+3^�g�h���t`���]��2�ּP�}�2G���r����.�:��S$㞕*V4�/�>+R�pW��n�����Ѱ�y��ɯ7�ŜV�(�#�hݓ^��ɖ�GFNH�SwFp\��f�w�[S���ƀ�RK�G#�~����Ko<���[hݜW���qu��E������|d��ɂ\�0An+���{�|�1�'YK�j�ZZ/��P8����[�C�}Mzσ�P����bq��W�k������Z�������s��>��K�
�5i�ߴ""c\q^�}2-�1���{~��,}H���BJ�[|)���3s����z�� ��l�t��]�7)��8�޽��z�k� �:s��[��Nk��������p� ��e�ԡ�yE}�c��|0�Y�د��0x�UעtO-Ո��g�Q����H��� zWl&�8*Et6>2�67�./dT�����z�ő����P1z�'T�P�<�v�}kټY��.�_�5��[m}��3�\I��4�R\0{��''��Mֽ��'za��;���v�8��E!�����S8`I���w�+��c#h���+��jO�-���3Q���]���P�y�)nw��ꩨ[�y0
�Ux~�̥���g����[�;��H��K�n$`:u5-�1�C�t���2�	������A���w�a#�W	c��s��8>����J1����p���dŮ6�n>�j��`H�=gZH��]x?皟v�;�¦�7��,�������֫�:�'�JV�~}{���sey�U��cѹ4�S����
�Z@X��I����>�ہ�QPۯ$7N��Q��)�#JTd��en� �,H^�y���V�3ހ%�{G�>�֟� ���B���<��*H�(���}��@�S~ooʐ�y� =�ѹ�=j6S�J~s��L#~	�La��1�M�F�;ԛs������g� +��<T&-ϸ�V��y�����\�Ӟ� )��zڕm�O�
� cg�sOT݃�����wt�;�m +L�v���#9���)_��1�SZ=�<S]���v�q��W���J����@�䄎}�R˟j�������<d B�m������z
��t��~�d{rzP�2L�c��b�:+ 	Ȧ���x���F�տ�fA���JTt���$���?:C;���G��^æ��FkƼ���z�=/H� 9@ƿc��V{�-J�)�P�}��X7ָ�YvG4R����̯�J��9��k��~� W���w��y �Ҿ~����_��� �|'�:/�mf1���O����ʹ��׊xV�Yj�3aA=�If��~�s�W�j��V�љG�Z7�.q��<]9`K�:
���ơ�8�C �9�x��ͯ���G&_��jԓ!ţA�m�3Gs�
���D��,�+�</�=KZ�Qk}��_J��;������C�Jʡ�;���BWT�t`�~��_
<7/�����q^W�o�ZǇ丹�F�Č׫��L:k$.�d#���Tt�������I~dS)9��V�kdpSn3�>ՙ�[B��dP��<�2>p1�a�xa<#���t�p[9ɨ�o�s�����%��ճ^��|>��� O�^c�+ľ�Y��s޽7��� a�F	Z�J�1Z�������
���uZ��ͽ�ps�<�^]�i��L�JH�q�3�F� ���1�����W�Z���{t�h������@8os^�6�,p�'5�6���Ӧ����k�O��c�z�9�W�R�]�ug�^7�O>�c�My��d�3�?
�~3E���8�!Г��R5���1�Z�R:��lu�4�VpN��_1�ƅV�r�?Λ7Ʃ.!+���޻(ғ��R/S���}Ʃ�po����[��	�2��yƫ�5'�g����t�leQ9ݚ�aA�T�#^m%4�jذ8g�׭��a����_\x�^�EB� ?GOҽ�\�e��&9��i�Z�Q�7\(R}Oj�Ջ���Bz�5Wy�uL�d����wm�R"e�&�L(әv�z���䜞���QJ��]��C����U�_�-�ʹ�xsRQ�\2��#�~����V��Q�V��!f�۱��;zWа5�����:�کG��r	=�l��� ^�kR��q����4��6>��1�?\�srsҽ�h���$�W	�[�Ѻ��ֆM�g����O��j��z����Wco, y��s��+|�z��2G@�S��<�Rq��²4+���Uo's�t�L�s���Y�=�ihV��z�XB�c�1Ld`��MY�+s�
`9�6zH����PȬy{zSU_#���@v+ Ϯ*ݫ#"�J���ۭMl����~a�Tq�f9��;��v{��{RAX��)E�v�)3׃K�z@�z`g�UB3��9��sS�<��S��>�f��m�������Vl�NhEe9��EUGniѳ��L� +R�h9�I���ny5"���4�z��������{�$n���C��:�ax�MU�>�3����8<
@?�$t����Nf��I��`"���Y@?/ӽ8?�לu�v�4�A҂7`�¦ES��-��$ 	�&߻�S���A'ګI9��!���,a���_�?�c�x��N݃9=�{��%q��kí��-�[p�{Ҭm�?Μ���t��� }h�?�E0�c������	������|����^�G��!��<��þ6��v��=� m����>���rFV=�~4L-��r+��W����qb���d.�Ӷ��*	*�:�
��M�����Ws� ���-��㪡���F�v�d�TN�Ҝ��zO�~'I�4u����+��ק���1OB++O�y��Kt�A�҄���cд��Z��>Q�m���?Ωx��%���\j��hxQ��ʹ�
r��Qp�8����{7�Gq]�m��+�ԏ/�Kg}5����LU�7D)�F���~��+D���+�����2#�}r9� _^�ǚ��Mz���W�wF�굏G���r�Ϯ��U���X�q�?μ��j��z�Ƒ�K�$�?�f��,KGQy���
W�bz Z�I��Ø���w��?����15j�A��e�X���>�ͳ�2�>�g5�e���"�A�$��緗�+��ԺM�8F9��S�T��r[����ڢ �L֕�����6�ǥq��ـ_�y*LB9#��ccK�V{�����w>|vpF�}�Q���|}�;G�4���\I�h���u+�C��j����1����h��]J74�XMp�:j�0Ja�����FM�n;��9�PY7oΘ�m��[$��[
H>�Vl�%+��G���}.ckx��NkDƼ�Y��
�w��̬u��-[�qg8�s\�����C�^�E�;j�npsڳrOcU��u*��~���'�����ڡu(�ߥb�F�E��Hrzf��F�9�*���l����qPqYKR�*e�o�J";H''ޙ{H��ε b�ӑҠ���g��#��X�8�p��� $��f�zU8bvo�\����A���S&o��t�� P��� z����m�<Uxs�S3`qހ(M˰x��,
6���~F�e��v�2h�֞�mݱ@�#�4����4�S�ޚ˞zqc�ڌnnM 0t�jX� �#F1J�~4����Q�y�<Ӹe���ր+37��szc*vi�$�犈�2 
I���e�������֐�)#<�ӕ���L�.Jq=����ث)�>���s�HD�60XqN��̋�t4�Gs�G"�3588�<}j��[�i&�=�I'
�/z�I�c'��2L�Q�P��/'��&�ڒC��sӭQ�G��O�j5��=@�{ׂ�_-W�z��M-O���W��>�2�r�^ե�[�ּ<F�KT?�$s�5��H��y��ןs��f,�T�F�u�B3� i6c�3���$��_D~�Rl��+���9�~�����F`�{z��]��%�P�P���)_J�|s�U����T��qY�֞��+t��� Ռ�6+��f����T�5� ��KV;�֚����-2%9�jF���我Wr��K	皈ꃷ�(�wJ�<5�U�N>��xzV�˹�K�рu ��<�� k���5��~�0����r���� ��ˆU�̬�X�j&�S<��X/l
A������׋�m
� �*��?e�_�6;���N�q�N:S�/�y�WRL�V6|� tU��Ch"�v�&������-��d\�^�k��, =�E����G;��>Y���I��l�dQ�� �Ul�֒hdV�+_Y�����ګzm���^�5�����c�{�s������il9S�x��1��Ns^��o�zE�����8�8�^*�Cm���[tqɷ��>OV͆� rz���>Y���
��sK��~FA�a�Z<��F��Z3�m5�֝�Ҙ�j
CY�cӭD��S���I�O�g#x�I��ǵG"�<T�F�C&6�$疧D_c6�
���%fV�Z�"��Ux����\2Vz��dZd���aP,���x�*��+�4/x6!�Y*9�v��<�*�F��Z�M�n g򬤬h������	�3�j8ݏ̽�J�H�995�B�`�sPɷ��*v���B�`I�V1�R�?)�H�b8���j �5�1N9�y`w�# ��1�S� 4���3u�	7zQҙ�T�M F���N�)��w\T�p9� +g����Ni������ ���*Nv������O>ƀ�����G44�n:����� ���i�s�ңf2>��Aɠ��ˎ:��9U���J`�e��J�L�h�je`Ǟ)���x�ښ��Ջq�i�w�?`f��S \/A��9�j�x�}F*#|
�v0x��s�z|n[����`�ژH��t/^���FqB���H��'����>�B��Z�����χd���z�=5w[/^���Ŀx�(�O����ӊ�@v��t���Ί�U��ǽ��E�U�2T�}x��! �N+���(̄� v�����}�~����X��vzd�z����ކ�� �^�����8���Ҫ�/�H8 f��$c����-g#Z[�X��8椾Ȍ�TZk|�9��3ҧ���m��c�j�;A��Y6|V�1�ӎ����%��k�?���}b�MJ!,��Bx�_�g�1�Ն+�>k��6����ּ�Q�a~��O�&���i�Hv�7�3^G�
=!���!9*�1�_!i����困��j���Ɵ��w_L��
S�ޠ���:��m��9r#z���� ~(K�M"E)\�!�^�{n�ͅ�ڐ9����|��M��֥�3����uɕ4g�!󋉛=zՏ�H��;f���CR��;`���g;1pGFڤ��l�� 9�_��[A&#5��+���x5k��$����W�Ȕ)��0���o��X����1�z溽jݗM�׎MqѶ���^�'���Z�:�r�@j����W��Dǯ�j�d9�Zu.7�5H�J���ᱎ���rj�^���ڑ�Wʔw��=oƤ�=�㩤a���� :Tdn^���j�!���j��O��C"�y�y1)�B��G���Ϋ��4��5�#�,�"ez�z�$�c֧0��ڡh�Ǹ�d�z�ZLi4����Z��0ƪ��cұ�3�¶�EMs#�~�����8'q:��3ڤRs��x�ўjmُ�t�4,�S[�f�\��wc�hhXtsҧl/�F�w=��jq ;�韖�O$���x�79�zS��H�i���m\�~4��#�~t�fͬsN�́O$}EFF(�6s�~�Вid��W�� �ʔ(U4��O���<
 b��y����?Zw��0� \����;G��X���iUS��P
K'���S�A�j=�`>�>��r������� �Ɨ�٥��^i ����#8S֞��⛴*����)�C7�8�}ߡ�v� ���L���FO�du�:�0�۞��:������Nz�ӌ�g�zS��)�Z�2)� �q*8�5�0���f���R���㚗�#�>�f^9��O�e^:
�φ��GJ��-O����|G�Gb���''a��5��m����\渍�U���v����Ҋ ����,�����F�5�w����}O~k��7���x�$H��<SNA�O�_Ң���u�z-i�l���¹��_iw[�u�w���BJ�4�VijЁ��.mltris��t�a�ۮsު��@��d�p1߁^��v�9��� ��_���n-��HG�YJZ�֜5<�O/$����zWW��f���G���W[��M�ı�j�,�^�I�����52*�B�j���S��ϋ��-��C"�`pEi#��J��u�4����� ������]џr��A�l��V��Gb����b�1[Zo�>� L�޼�R}g
յ=KOա����s�]���!��(J���k�Y<L�am�9���d}kƕ.���=�S��e:���x'���կ@��Oz�u��s�.�b{�X�8��sJ�w2n�b��*/+��Җ;m���5r��h�+Ql͸�jΓx��a�����-�/!HJ��46�ޣȠ�=���KWV4.�\��,��y�2+"=Ug�,�f>�W՟��.�(�ʧ��_E|'���O�Z���+[-&ь}+�8����e&~w���w;�0x_P��FL�	<z��9��D��ׂ�0��A��?�~�]��̖����UB ��_�?�ǀ|!��}6�%��� O�WC��C����mf%�֎r1�����T� T�m�2kԃ�<ʫQz����ޤ��:ՙ!������L�TE�֥���9��7v�\a�a+�x%'��+) ���E�p9�����.٧7_N9�΍�*�=z篥3n�$��SDx�+tD�o�H��qRyg�g���� �R�'�b��}jʾx���c?�S�,=qVc`T��4�7��	z��_CGO�
~N���,Es���Jc � :<����B�Ҙ��S�6܎y�L�on9��t�A�������q��&��.܁�=j���@?��䞟�+7#�b�[Qe�Fi�jc�� ;s@�|���P����X� ĩ������z �d���Ҋg�c�����3Q���چ�{SW�s@C�y���6�H$t��l�8=��e��@��ˑ�Q4g�o�y�L���>��P��ӕIo��@�"�*:(�+'S֞s�2���C��(H��x���ӊ�,�TR+�s�� V����B��'��f��ʖQ�ǥ U�N�)�W�2�w�ޮc��	)�]s�� &���#���A���� z Al���9��Q����+8���fM�߅'�G��7����{՜�,F8�dX�RG5��w�-��A��w���I���l۱�Hw/S�׊����\h�y��E0�w� O�,��Aߠ��-��׊�G����'�d�Ҿm�
 ;W�x?��ܖJ�N�3�Q?�v��G��#�F�wz���K�Շ��j��]R���R>Ӟ���N�Eߊ������ {��k��#����%�V6��:�ƷP7�����@p�߇� _�zcK8��� �y_ū�][��� ���f})�_xf(|�T��[�M�O�h������G֮ˢ	�'���<�*�)�o��9>��*n�5mlyO���� ��O���8��1AۃZ�f�<M;)Kc��X�&����ᶧ%]��1�k:}�b�
��ˁ�j95`�rsS(Ŏ���&�*�sU汗�+S�T73P�0e,N@�{V����՟S*����Tz��e�'�O%�v����I���'&���W=r�E�fݻMh[\c�c�CX��U���_�5'��X�j�(Pz���=���ڪM�Ө�O�}�V�=��#?�n{g�<Iyk��/��I+�ٯ��Ԟv�co!�πc>-�Kl�q��3@������0U���4RV>����Y-��t.�\����>+j�:ż�I)����ֶ��dۙ�3���!yo����6�tӍ�9d�󽎛my�K%�|�?)�ՍoL���Z���{���A�J����VZgt�٣���܄���O4sHݹ�]"�4�]�=�=x��e&k6Y�2y�\c���7V'��E d�OJ�GLRD/�� j#��I�_�9>��z�f��tD�ٙ�aijq�l{�zq���#b3�� �jh�n{�zTJ1ޞ���5�#h�d*ʄt�G֗��?�Ԋ ��e��_z�ŏ\�n�ڙ�tے=��3|ē��� J^ >���2��)��6`���sٺ�e��?\
@P�aF�,zsT�H��5�^�-�{��.�a�Ҿ��W�\[��kY$�(ɮy��v4��9�Tf>���[���d8��+�cM�S�Y�/5�^�Dco��s~5�}���yVxw��1Ǐ����4�g�B�cc����eh������^0Ӭ�ۧ�{��p��0�T%�c%a�#1�֬�K(��5I����4�gېp3ҵ$�۱�}�$�6q�i�v��ޘI��RR˷�NPW�֢e9Sч^8��s/�r(����2I:��9!� ��$V�L��O�+9o�LWّޝ�=N =s�w���� L��B0��x����M�Z��|�����Ὠ h��Ǩ���Tm����Ym��P�� �� 1�<���s�����nڹn[�1��NzR ��qMQ�H�Zz�U�M "�v��$��Zv�'�2�x�P�]��l�b�Ca^�a��_\W��d��d䜟ʽv�TU�t �^&�ǯGcL�>��0���9��R��%�|d�luX�0nM	��x<{�OAY�~�����昗��+��Bх��u *��!��ҿI��<W�<����Lli擽w����RX���wz�K�,�e-��5�ȤP�jZ��|`�� 1��#my~��I}pd|�}i>o_«�|��fұ�97!,�VL����EՍ�H�`�s�~7��t�{qGB���澒���!��jCgou̬ќc#�µ��#�8�P���ȵkX-��s!�H杠x&�Ĭ�I�j���Z��V�F��#�D�d��?���OGk[�FŒ�#~�q\5�{3������ �����+ָ���VJ�Q,�%�ܜp 浾:~ĺo�/m�B��ة�ܧ��4���'��m��Xmp��c�jO�ɠ��O�ki�>��H"�޼yW���:qzX�A���GI���3�k�մ�ۘu��~4���� �]�s��򯎼yy��1�Ҏw=�k�8R8�+F�y#"��S�=�Z�vdq�"��e]�?\w�^՗M�R�� �N+6@Ăzb�ƆI��'�;_@��>��~;�e��W�]���5u�~��5�6�u�%�TR-���tG.�7���n��l$`����x���K�ZERW=Z�k]Pƹi�j�յ��m���m
2��'V^�GR�����Z��Pn��o�'�G|֊��W�MYUi]���(�8��+C/^�i�y�?��q��s�z�R6�u�TR.V������_C��W<���q����Mrv�]�w"�����μ��w �x���9��I����=����T{�du�c`�rr�C�:������:>8#�1U#�wXY�'��a�e�� �+.dh^��c g53;z��Q��ɐ��1.<�*�[ل$�3�=j5br�ڪ������RCp�H#֤}R�O�I�y�^���X��B�����J�/�G� ���PN8�gMOVk3ޓ�u䄖���վ,�_+�M��+ȍ���!�����^*�Q�e��[Z���dgv��}+����3g֬<�Wq�Ugig�'�����Eha&�Z]��^���p8�U�E���Jw�� �y�T��'<g�F�P;�1Y�}�{b��(c�)�.�c'����t<b����ŏʧ�U)�LI#m�r�����
J��?��L{�������6��#�Ҁ-��{���"ƥ����\/ʪqCI��ր'�@��Ѵt��o=I�}�v�:sN[�=�?��e������ �OS�9�A5��������OZi�����j9� ���V:��Fv�ҝ6������.ye�8�{�l0���Y5%�r>�Ϸ��s�cH,���EV�:�Q����9�J�oy��H�E0"bW ��ƛ�3��l�n/A���Ua�����ÿ�]N�Ú�[ȻI�z��[���xv�ˌ;)�ں��#E�^k˫fz4�⍯�I_h�H�P<D��85��<�{�WJ�t6r�ݻ�b���u����ԭ��&�x�Um;X������A�"�_Wb��=K���6��?��|�8�+��7+m.BH��c]��Z��'��񸯈�����i��N �h���I��@U��Uo>daڭ.}*��� ��Q-�i|Clp��V�>h}*��ܞI�W��Ȥ�._B��g�Z��/�dZ�%k�U�h�U�����ӵ(�A�S��"�� �� .��+m�b����������Z��z������My�͏S���g�_�����B�ֽY~:=ׇ��2�x��|�$q&�Z6�q�s1��u����}�����$��k�;���@#9n�� ��P�+��A�����h�.��o�|��,��'��y�)��9ݫ$p�5av㞄����&${չ�5�#d!�.��ߪ�j������wA�jz���r%������pJ�)U�zW_�/�K2}+�F�J�)�yܼ یVu�|��ÖZ��t� }+���=˖G��U{�<w���J�la?�f�㯥5���:��*G�z*k6nI�6^sL=�)D��t��%�?�O�S&a���XH�W��-����i3��z���+	�Mpq�K�)���5,h����+
�t�������d��>�@� ����5��gTH�̉��/J���zXt��lZ|e0��*Ƚ�zgqPs��YM4���|��)�Sd����r�MntI+�U��#�&N~QY�:�z����H���k+T�n�j֜�1�]!��r� �ub{��y�7=�)<��̄,Mv�
���K�t�����Ζ�e����\w:���۸B�t�J��\�mV튷�k ö.Nz�]��<��cvth[�E�I@
��5.��¶���ZURPI�8����i��r=*�{�T���]����)������Z�W�n�ç8�I�yq� ޹5��bV����`�O�
��*�DS�����m����<��#<���ʞĕ��oQZ2��=+*$i$FNkz}&_���ӥ$3�f�#����� �<b��/˃N��8�%p5�/�Y2���T��y��6��~ݥ�n�X5��i2R:S��+���@c����n#8��+���������<t���5��&��ڼqe}����Y~tt��$[������zi��jŤ�q˜���Y���]���@��!����ێ*�rr9����*Ȼ��5Iax�+�k���q����Ӛk�;s��j��� ��#��m���t�a$��"��)Cpz��}�n��\����Z0�W��Z^��Q�Z��v��.;�&��h��E��b���'�H'��u/���.d��q������eH�=}+T�Ե6�-b�!̇9�c��^��0��3ּ����u��8V\`�z���R�A8]�W��t�
��<�C�F��I�ڊ���?P�#�(�sۿh8������|��y<� Z�����v���y��"ǘ��}�h�1! Tf��o�v�x�=h-M���Y*��QVR��ZR�ڟ�2�����#�ER���==�����Jع|ev����hIr�����Ȏd��T�E<A]�z��B�A�.er���v���޺ox�4uQ����E��nO�T2�I����:��Mκ5aM�3�����Z�%Ր�8�k��-�8f5�Cm$lIc���f� |��W��:���E���yc������u'?�yo��g��v���.ݲ>ls���b�ϕ�q:\���3RW��9�㯵T󼱷�s�_�R4%e��Z~�>����±���V4����:�qWY��=7[Tm4 A8�,�:T��R�F8Zb�ߥ{�H�%�j�;����95z6*���W� }MoЈ|E�=YabGNjc����b�Xl9?_�Z-�e�t����T�~cM�@!��������5`矦j-c�g�X��ڝ��V��fb �>e��z��l��v�?L���x<�S����U�1��ПN(y>��F^;z�v�|f�h�n>oҜ�#�����mf�8#�gФQ�?��8���~�Ky2B�?�^b˛�0I��}��>ƶvp3` �ڸk��uM;}8�#�+ϵ*q7�6���7Pjl�/\��F
��J��7^g�X�)�ri�֓X�'�6����ё�+R��D2��\V�1����^.�c�v�����?N��x��T$���\�(O w����U��a��@�}�=��������;s^���|Y�9�k	�r}B�nLx���k=lda�n{v���ϩ�֨�i&��z�Ɨd�G�U�̛���g�t7v�,X!�@�PY���MkIj���9�#�3�<��Ԥ�RV�eI��o��zÀG&���>ܐpX`����AJ[��B1���n���k�c��{me�m�T�SO�D>j/=sN�hO��at-dR/�+^}y���8<� ��e��L�����ݫ�Դ�-��G.yf�?#q6�^m@����*��Ӛ��� R{T6Y�o�@�A#�Z�����)t��"[�1�9��J��*�s���I;Cs���H��T�ӁQ�Lͻ�·�7f�+3|�9�
.�ކJi�R�*���#Cy
�dc���{��I�1��;U�	!֠# cޯ��c���wu�zҳ�$�,j�����R�D��^\c;�v��|t&i�4�=>��R�ʔ�8�u��"@sYWWM<���x��(n�Ƽ��s+n�H1�ӊn,Q�d�����X犻>�pc��I��o�jظ�e_֬��O�(O��� c�MA��\���ס|1�Ŝ��`Q\�ed"��Dwu�$�Q�zƠ��*1O��<�ګ�:�;{v�oa���;4�+ֳ56�D����3�kk�֮�AS��� �ꇆ�n"�<q:��ps�hdy�ÛP�����e'�{�j�׋����QRƏJ��>kc��W��唁�_S~��)�by$b�X� ����a>��|D��Si�{�4�}��
>��JZ ��{����8���
�4���?���岣�J�{�C��S���Wn��'�Jع|f]�<�kXd :�ɋ�p�e���DEXn��!��@$�����?�e��#�Ԍӓ�Fp�1��Z]�ȵ�����}>��Qg'��ߊ�k�hw_g1����+�_��<}�3�Uk>e��˭��e�u��u�ʚ����We3�5�k|T�qg�TJ�?��%���Ӄ�s�]
v�|�� ��p�SN�8����h𮨽l������4��R�����░�'OF� t�+��s�t>ao
j�Xa�����Ï�I��m�.�s�_,� :�FO��D9��*?�G� �K��a8�i��흶<RN����*��ڙ�l�$t�{���r,T� �j�?�a��x8Q�ꊲ9$��c�����c�>w�6��Z��ukTKaqc�Ȅ
�:��>��+
٪n=�+cŚƛ�xfg��Hd#s(�ӿBcd�|�����0{տ�Mh�+��F r �`�k�;�>&&�M#�J{!��ƙ#I��F��e4�~\��L��e���?��*�ӊF_j��;2��v��3P�gҴ���#4�+�~՗�6�R��W�<B6��u����+�9ڼT�F��1J4�o�py�5��-�Y��������G�G�&H\�]�ڲ}�B�F1^mjr����U�tl۱���|�I9���?�U�����(��yM��%���MzXC*cʩK�:}�e�=��B5d���G-��ڹg��5�O�.,d����ku�)\H����^i�rL�u��"[��#��K{�7dG�����uծ�$�U�!S+х$�8�W���o��G�c�:+-���خ
��S�)8�8����X�Q���V��Ө�s�`��>V�i<y��c�W��x�f`[p_A�nG�)&�W8S���s6���佶�b	���kQ�[�+�5溶��r9o�f�Y��{U(�z�f�F�عԐ�[����f���<;yyn،u�sU��Եh�A���z�\ci0�� v�#�]Q��s�\��h���/Q~�".~�
�A
i6	(c�+��'�h�-��E5�|Q�nVqr�q�3G�����=A��c��T�|�;I ��s:F�}�L���6z*潒��:�ǇH6��B�]r?*nnZ�?OK�Q�]7�|45K�XeG�Y׾��MďqnQ�쁟º/Y��1�1Dh�f��u���xb������=r���p�����f�OxC^��Ie�r��Y��:K���8��5~����4|�y�Ia3F�N;W_��}T���;���5����+��W��6���)�+	Ժ�9{�z��3Enϸ�{V�<}�i�Ks�y��]u��X�@W[���46l��r=E/g�����ڥѶ�/�ር?�]k�D�@�:���4��u���$���]�� k�B�-��3�JӒ�9]~6��ً7��\}�af��f���b�,FN3��y�����w�qڟ"{��z}��wQG����Oi" ����
������Z�	�mX�����z>���X��UB��W�\���wc竨��q��O�j�9����	�hf�=����.]T�ڹjS�DvӨ��zu��o�$
ӇV��2��&�r;�bQ�=3S� j\m<��5��coi�t� Zۜ�R=sV�o[jZ{��Ň�^�(l�1�kn�_h�!�<V��7��U"���_�Y<C12��{QP~��Mu�L�p6�򢲔\]�#+�����ē�d~5����oc_U~���dq���𯕷~���{XO�6+�F���$�����̑�qֽ��� 
�K�u��cչ8�]���nx���?:rȬ3��>��߀�v�w�n��G���M��d
2Ts��R��ӱ�K��k��߯b��.FZBq��^�����G{����3қ�������?Jк�p1N�4��ks��uO��xZ\��m�#s{R�h��r�ʾg�jGplW�^�3�M*�1�4o#�!����~
�cP�e�����J6G�Y���R*Z�.H۹^x��൸�����^=���RKf�������QI�r��N@�
ҧ�gMY����MCŐY������k�O�� �JO���1�S�i�,^bZ���d�x?�.����}��n��$��^ ��/��L��c�~P������=�%ȴ>���6j��I���+\�!Gf�G~;V��_�Z<>f�RHyc9���k���>$��K�UD�6wנ?��9��[x�X��rF����%c����"[�6�<��1�x�7���E� ���{�� ��t� *����y�ry�Z~���ug���x� �~�ϔ�t��<R��r\�?l�/v����f)�����O?�zƥ��K�v.�h�K������Ҽ�kI�<E
�A�T�0���c:�4�:�C��2�`�O�E�1l�^���b�>�Ե�#q>z���%���7d)�=�]�<yq��*D���N@ҳU�ܩS�C���C����~�*pZ1��k�l��~B:瞕w�'��֦��9�{	�������h��vy�4g��.�RP8���� �Rj,�>܁�?:I$�+Ўǝ?���s�J|1�&Dv�H��}��vZ�����=��/����:�9`�X.8�[�Ҕ��\`����Yi!�?r?��œr�9���Em�i�]�Qn+�!~��W�Z��S�>$1N<�7n\�i)\n(�2�9��� t�[�w
��+���>����6||�P���m<�9��a=	�Rrh\��M�ڹ`S؎��0���(�{_Ə�v7���Vl�  V��� hZN����K7�AK�j'�s�>$Rcԩ�5U!vp�������O Xǽ���S����R�ceyo�����A����N�VG���'H�Ɏ�U��f��\��9�v�i��wAы߈���|�ݜt�֯���ky"ã�����;O�*��1I����nd6�9�6rq�q޽��^>ӯ haӼ�Ap�n+ʧ�d��p��1RՄ�8�UkL���$;A�O�c<Q��1W��O��W�߼��q�JqcB�>�\�lf�'��k5���f��_J���"i�v.zU�%I��H<��S(+��̩�qZQ�Y:����g�nsY�)�MkI�;��#�	�aY1ٙ_b�O^k_Tb� �T�����JnƐ��.X�mN�p�g$v���Ě����&���*�8��{Y5�-c8i.G־�𮋡�>��\y+$젴�:q��9v;�����~'��3���s�x���Ś�ы;�<�^8~u��oŻ�Ǝh�,�>��|Q���j�+'������Ri���~���C�k�!>�W���B����ai�9�*���+9&�������}?�o�曧�_j�w ˬ� zg5�Z�=O(���k�f#g�a�=~�����i�AׂNs^���F�����FӍ���
$S��+XF��R��=�E��������_|V�Z��,1��<י�s��y|�9��*h�hGp�q#;A=�{��(�C�0F͟�}�b�z�m��0kڧ�v����ij�kes\�E�{;Y�~r� �W�����y�X6�p~\�סk�>���x�U�!T(?t�kM�nAa��Yr�shx|:�.�����J��ýz����4�S;� ^���6׬�X�,f���};���&��=)no�mv��H?��T�$8����ƍF.{H�r1�kɵ�y���:V�����U��t�;}Id�UE+��q�¼N4-��MJV=+�ƋoQ�F=�v��{� q�C�k�|�NA�F�S�C��*�C�I��K�Ǩ͛X�Ԋ�9"�>�j
�!�m������O�*�WR�*1F㺟$E�.�-3OhUc��#�jI72`�O��&�g����v�0��w�����X��2���s���Exu�6{ԯȏF���k\e�־T<Hry�&������f�����{��ק�����-�J���ÏZ�ˉ���-���^85�Zl��F��F}!��[k~�^6�u�������|Qv5O�^w�澈�c{��.\2��}����#A��3�q�rT���W��.�XکHX`��zVZI�=��cH�<G4��#y+��Z�;oG}�H ��ʅ���Ԟk�v$�9�a�wy,�C�w��J�+"b��'�3��v�;����(o�VuN�ן��A� 	ᛝ���-Ơ�
,�ٺ�����o����vh��I2](^U#�?
�=�إ�#vEqV�u��V�i����ȯU�k�Z7�P8�'r��������j`��/S[� �ƍ�p6��f��@� �i���F*xQ�n������H�6@�k��u�?�bLq�Z�>0+Z��]������`D0+î� N@���r��Q�UĲ_��	�Ԟ=f��X��W3�=v+��g���]���kK{PP����p�cvՌ�[��<���L��z_�nd  #�5�z'Ƥ�mDb(rx%������H�
m�1]1F:O�Z�˧H9*�y�#�c$���=O�,=����mn�����_��d�3\ޝ�x�'E� V0?�M���sR�4t9�������-�^x�V�%�?�@	 �<��ֿmm�� c�1Jlrfo�%o�B�p3Һ�"���&�Fa9ϵr�<�-56� �w��}=���ޛ���Zm�a��ҽ�)�=Y{�<�-5ip����*J$�c�Z�V��Nb�<�HН�޺ԭ�����=��
�bs�~���[R�=ZQ6��ks�M�w�H�7�޽�W��:�0����p����*e+1(������4�$�Z��AT>2q��.>����E��Y�HcP��ظ��<N����\l�O-�Ln遚�J�}�s��}�u(mm�1'�W�i�X�9�r�73��d�v��?��M�\�r;׋���R��+�b�k��������z d8���׬j�1�(1'fp�'����2]B-�.͎k쏇z~��e�H�	ʿ8�ކ�QV>j�ƕ�_x�Lp\2�܄�}�h�H�`K�������Ş�JZE���ּ���5I�U����^��w�'�+�S�$��М�� ��ڼ���?�3}�����n<�����	�SZԴ�q����ݟ�kTӵ�}P[�3L��W ��Z�P��#�|]��'�zl�6���܀Ex�nt��"a����O�>�I�s�~�����J�Clڤ��\�u�_c����Gt��%Oڜ����JM#���I��)�9� Q����A ) �U�#n�hQHxg�>;wh��p�3�u��֚��5�;�ޱ�K�V�(�A\\�9���Q�˦�#s[���kR��g�d�!󏹭[m�X�"�����Q��_J�a���sWu�=�튥d~l1�ޏ�\�u��\�y*���ױx���xeyUa���z�,k�Dd`S#�{ǈ�Y�`P�m�i#%���Ȍ̏�f�&��i0d9=Nk~O����-��yY��H�������M��u�+o��G������1�;��^�� ���L��P.<�`|=����KQr����x'����1���n=sQ86�+�����v�"h����ȯ�f�A# �������g����=����I<�ޞ���~\@�үZm�V�$L���+���{)V5��漙���S��G!����Q#h��˧�՜��N��rQ�I�6>����%vu�@�#�RsY��;��p�s~�Y[*�eq�jQ��rz.��U�ܯ��;�{ףxk�f��j1%����	���y� �t�t[ǂ6��$s[�4[�K_���F�Nx^*d��ί����]� P?�5��W�|^��-���k! r�x�xkf�LH
� �5ə@�i��{�j�l`0s���J}���v�Ґ�ޔ}����c�4�7{{��)��֦���s��D����LͶ:�[���7��^���C�߃EE�;�rc�v�G�Exu�6}���D�-�\�`�_+nď�\��_�,�2� �k�\׭zX?���{�,d�G#�l�5��B�d;_ng�x�8�J�HW�:u����ǡxo�&ܛ�k��'���h�n��6ׁ�=�e��T(s�gȓ�4������o�a��E~�#������4-?��Z��1�U�u��=�nW5zO^���n���k������eݵ����Ey����1�`���k�� ����i[ӭU���"�!��t)�x�2X��[H��大�� ֶ�|5�]*C��86N���f�\���C�GNzV�����{V9��%��&��^(� ����0ۻ�+�>�<�HFw��9��Rǭzß����O�\��D�I�7�� ��Q����RJ����j�g�w����J���^�{�@��*3�Ve�� ����#���}Y��#�l|#��Um�|��`�U�/x�R�Z�f�ֽa~6�������_���G���1���I��p��a!�^i��'�Dˑ��G�{�.�;�
�#��6�ݩ��5V/�'�A�w��.�"}[�e��ƚt�$v�Xu�^�� %����� �.��2���i�U�g-7��s>��r�w�,��� Z:�m�ֺ�5]�9�;��'ǻ��Yb�:A��h��깔a�C�;�� Dd��HS�z�>�|7�6[� �&Xz�&�k?��j�1rޠ;U|r��,�tl:*��B�#�O]O;֋I�I�g<�=큘�QV��k��C�44�� ����tb��-���c�
͆�x�ǃ^�E�Lg�Nj����x������8��S��5;�:�l�ݓ�}ӫrǁ�-�����K�|�qU�<a�7���l�p���P~"ݵn����������)����t!D�O��k:W�m�郃^,s5�c�k��n�<���i ��oP�ux��8���ʹKC������$#$��J���Z")`��s��[_��Z��z�r1�a��Q��2\B�\kk} �h䖆	6�g�����LȲ0B��^�}�Z�V�L1��GҦ��c�d�]gc܁�T�� �}�K�֔c���jF��{�)�&���H1��_B�s�7�c�Y����GQ�n��W�^~����ή��pqSi�����6����rł�҉Y�=N���Kk�f��*c ���1^#�����}�:uā�\
�U��-�f��=I�ʶJ����wڽ�^
�J�Ǻ4
YNsB�v'���*����~W�f���S������ò��z����b�[�G���п-�~Ha#�������o�������g�/� ^�_��(ۦLs��5���!)md�
�?�5$�Tn���mc�o���|5�L���t���t��T��  �s�z$?�mf
c��Q�Mu���ᕣ�/���ҹ\�G����9��o��@��j��O�H��q�>b�+�d��ȅ@C�6��w�o��r��Y��vǸ*��*wkc�d�;����+�T?�<Wk�=���Mz%���_M�uš�N�̈��=k&�����6�,jQ�?�S��k$sv?�_(����u�����-�Ɵ5���C�浾�c��u�b��s�W�ٽ�Ln�q�̟)��������ķ�5D�V�ðC1_�!�}x��/��(��܍��U�%�h�4q�34j8x��BO�V��.��U�n_#�ʐ��L�I��=kh �Sk2\�]�fj͗��]2CNұ��֕� ��gc	��+�h��V�cw�ZJZX�<����7��m�2Gs4F����Q��3|��3�i����	f$ƴ�~3�^@)�S�����@��Q��S��5����~/R\�XեrE�L����D�G��am�_�z�`,�{������I�I#���y����FA73.=>_�L��V���̅��'�̵M�>�����[�Ǩ<2��I�Q���j�v��l��n39���g��Vy&���2{v���m�I�fu�.����%��>w�TY�=�26�F:ױxO�E��f��e��]U�¯�z���������-so້�Eq�*�����\���u|r�^�0$7w� �א�^��>U=r+�m����9�<
�m�L�XW���qIZ�z������7y�t�n}�q��Ls��oxÞԛk�y���=����S�E���w��دG���?I�� B�"�c��^r�TZ�/��XN���w��r1�Rr>�Fd���M��{�b��S�)�N��c����u��wV��4Uo���d��7��V^�>����U��aۦ9��{q_)��9��k��l�k��3_$2����]�?���n+g�%8�_Jo��y�Ԙ攰��Z����c����S�SZ��`P�4���>$S�c�޴n9���T��1Wnq��ON�+cI�F\1퓯5�;G�e�m�w��|�J":��V�s�Z~����LĜn�e����h�7��k�D��88�&E5s)�g�L �߬l@�}?Z�?e��0﬑���Ďi��!�ZN���x��Rk���g���0�y1��X��5������v�������Y���)_�i��$�/�.}
���5�kRP�!��n?:�/|]��O�,����nN>�����*2�ug9 ���_jՏ�oIc�P��x�V�.&=�V-�#j��<�+���*��2L�$��m������U����YB� j���O�t���&�p���/Z�O���̈Zl�H��F.G�A�6ڴym['�Q�ˣ˸˪���v3Xme�;�[�Ea�V|��.�I�&�Ane���F҇$�搌�dz�3��k���?��o�uN�-�Z��B�E�\q�מ�x�����5[k�6~W�V\�ƽ�G�f�}�I�0	��{UA�&�$��ූo��4LrV�,kC\�˩LH��T$��z�OC���/��@!_�F7~��ĭWJռ�.d2�P�z������J�劓R���>,XE���/5L��,3��Yr�z4c��g+���Kq=����wy���<瞘�����L��u��y��~��#_�=��;;Ht�8�x�n?���"�lmuI����H� |��׊��n�>P�¿��>�"�4k+�����w�t���_�߳��� �:Z^����hf�$bG ��ү�����Qso{1/4�F8��?��Oi�Xi�?��Ձ8�SUN��-��F���W��3�q$�n����� �^C�W���'v�[��.(a's�ƽ3��ǇIH��^qq���J[�Eܯ�8��94�s�Z����.�[�x$�S�����>��h�-��NP��W���u�Oi\�U��6gڽ��Z�u;�k{M>��7,c���UH��Ѓ��V�y�����;�*�w�'�S�e��<b��-e��a� �6G��~����_~η7�����-4�_~6�_�_�PO�S���� �iZوh��s�MiN��;0�0��� �ֹ��3\��5��
�U��\<�:� ��?Z��I�O��<F�qW�����wc�S��O��C��/�B� �}�#�c����� ��N��,e�9�]���7���t;�z�ɻ�lzr?Z���o�u燮r��x�^���}�$��ߝyk8�C�Qm�5i?g�����2I��5��xt:�kf�kꯆ:���ʭ�x�"����?x�3t��%�s��B��ԧMX�xkk9����EH�ឦ����?��z����㉖�ʉ����Z�¿����V-�zM�'��u:�cd�<�E��}��,�F���'�ֽ�º�֭��h� Ae9����	ۥ���Jʬe �|dת|�2/���#��Z�u��b�(�����z��<T����&V�=����4_ه�G�_��kҢ�u�!L�`���3_7��5��n�\�pⲾ#|NՏ��-��i�g
���˔TU�����,�+���؍��%%#H�?�{^���-һ���`H���<yq�$Vg,� ����.�g}%��6Əo-ҽ���VwzI�
���⍵�쌶�0Yx��}�o�����l��,��'�?y7}ޤ�����O�|BY�������{ŗĩ/48`�]�'+�k��Gc��Q�n�7�<A�Ʋ�'�+�zVϏ�Ԥ�[�Ydu+��`V������c�ٳ�ڷ�/�}���.6��A�\��F��(������H���0�9J9�4�dyCu���^��?xz�K2=�^�J�id,��d���M��,|ǗK�2��GZ�X�r���9�.��g�x����K�4�-��٧n>eo�z}���-����H���� ~����R�	oa�J�m�0�Yԫ)"�ӌY��|/��������ng W�߱�����;����O���W1�(��	����:]�
����j��ύ%���qHT�)�Ohލ��*�O��M�T3<Z�gk�b6�0�����_�̚s�2�c����Ck�:����$��5���K����'��~�q�W�G�8��{�č�Ы��O�:Ey�>x��;]M��'��i8��w�V�,z�0�8��� �����Ue�;�(9��W����Њ{�����G�i��l�����#�b���ه��̺L�D��8� ���%�4{�;{m���P1��_���xR�����I��o[����{����G���KS���,��I|����:������%�R᳐N5���R�R��7��Q�0�4���\b�V�/�W¤4ҳ:u5�BS��EXG��w�Eê�]����/���X�U�S���+���j�2�:��j�����H�5��1��_��'�(��_
�r,&nÊ�|��ٓ�IZ�|D�����
�N1��~#'�������;��D�4xƟw�.!h��R�2{��^��I���@�C^T�<���j�ф���F�65�q�0��|������G����+ȯ�ܥ�#�>?4ܷ��+��D�G9��� h]��M���ۃ_"1>c��8���qc>!�6������W����'�Eo��5s��{�^�C�� �JFy���;#��x��2�.~����5"�F�e弐�O�W�h�  ]Ce�Q�ݴ��Oh���#:E��!�r+f�5qV��7z�=�W�Co>џ�WK��;��|D�Q�@�`�ƾ���t�Fd�<����S���:��8^�c�U����H<��/�V�A�I�� -�V�ß�x�R�nc����8�v�����w�ε�(��h6�fj��~��G�ig� (���j׼YØ-��53�}�]O��!i�6�ky���+�s���/ib�#�6WS��S�1^��l�
�I���uf����(;V���ծ���:V���̔Z��P]x��	��EԷҾ��;��!>��M����>���=��� �)Ǹ�j�g�$�<bR���RqڼLT��=�+�D?t�*��-��j��,V�4q��|\��v�0�X�ے���t����[�:�k��� `�g-ΎX�+�X����?�^�'�3���I� _�fA�pz���{�>�h�-�ͅ��o�Z���+4hp⺕iD��L���¾8[��n,� ���r�j���='X��Q���B�UR~���i5V�:|
���r��Z���?�:_����V�2�f@G_�)V���"��ľ���r�N�k�d]7����U���u+�`��҆T���;���xЌn�׊���h��� �%	��1�逸*���~�|#�5��E��{g)7�������M�E�2����|c�%�/��f��Ant�x���`+��^��<�G�x׈v�1�>n���9�.�b���gHzר����=��~�������-�Y��M��R�x*�������e?z�~1 �b��Y��G�x�$� �1ۺ��;��� ��l.�C1n�g��>����.�JF�'����U�I��s/����_=$�{
�Z���[V��+���_:|B���j^u�,�f}k��
H������^9�m.fͤ����]wiX�y� �]C��ch��I����HO�^���/�Y ��-^c�X�~-�n#^��Վ(�|��W�;�%-�B�:�_A\�l]!R�i���9����v��1���y�x�y{瞛My�V=۩�v��d����[[�:�\`7�7Ə]x�Yi�f3)��a�x�F�C�ƹ?�_i�H+מ�ׇ���z�h�r�[���*�
��n�D���·�j�q	�B���)� �?�w�=�o�p�6|�����I��V���g���ֽ6��Q�a�d���o�ǨLK����������7��Z�*���z�Ҟ ���c9�T<Hѷ��i�U�����k�M?O��g�$/�sVO��)Y[��9��S���c2ܴ=�K�k�Q�Q��p+�U�����䁚�����M�p��^Z�F���,$���чnkK���VV�Q[������U�����v2:�'�=+��W��=Z��,�٘cs ��U߆�*����I�H؎y��"�{�s����~>S6�(F��r�/��W��ywFz�+{�*K�WS�8֔a���"����m�Pc��v>���5���#RH�����ulx�z�ie�����sF���B���{2[��Sq�7��v:M���Q���+���t-�U#� ���ȦZ�T��N�S^V"���7�� w�&�r��}+���yǆ-UW)��=x�𿌭�5�y�	l�?�w�8���������FF�\J.�E���9բ�G����^B~iXs��T��/st�L<��� ׆�[��#��oR��Eu6?�YG6y?�h���^�|c����E�\�c;ca��W�����p�Y%��V<�t�~����*$���rPx��^�D.�[�8ʠ��[X��CjW�� d���sY6w1�!/�ڲ<E�J�D&)VIB��"���4wT�PjcN�sF���WS� ��v_	~�&���c<ׇ���o�\F�<�p:���:�q���ҽzj�8k;�GĢ��al0�V7����*>�9�?��3�T9��+��� �\�]�w`JƷ�^s��ơ�3e��k�4���J^I
��母��r��I{�a�X�ʪ$��c^tS=F�G��m��{����-��z�n+��?�$�`�/�u�t�&��R�|�.���p��~"P�fݑ����yU��B����k�[A����]�Ï�x.�3y*���\���Y6���2���#T���^]	V8x��6�����_��� �Rϧb@�#oZ����C�E�� ��y�_�g�K�@N��j�����ݫ[Ɔ�q�O4�[Vkr��MR�h���ו�>�Rꚵƭrev��Z��N>��ec�m6w�$�u�wd0�4S>���R9X�𢼊� =�=���Tm.C�9�+��d�~c������%�lu�����A��ƺ�ǋ��mX��s^�i�jo��H�3���J���Iu3־��sw>��<�j���+�{�G�� ��]ꮰiӀϞc<s^��7�|6~��d)�s�
��	�*��T���"�HR@���Z|�Zy��3
��ˬo��ͤ����x�[=bY�;]���5�~ծ<Ad�M&X/�׽|ر�O)U���7*M}�GԿ��ʹ��B)�J����~$0_N��?:��e{5�����a��h���N�_�il�X���W�D����m��T~��>���to�h�����p��՝�?��/�`{�:�IFK3��q�m�ɡ�M29%���֪|5��Mu	�����x>f~j�ƍ�p� ��홡�m�X����[� Y���3����cj���Âsֶ>XOr�C�\��+�˔�=F�Tվ��h�m�H���Zx��-"Wf�o�+������L�u���m�����  $W������h��;��5椃9|�^���B�~G~�����1��MԄ�G�s��]��>6��+ۄ�ˁ�J��7s��'��/�]斫�qF�r��?Z�5O���pi W���־-���y��'٤tF9�I�k�U�3Js�Ѫ�"�O�n4�R��K+i�ޱ�U��f�:�K��_��1��w)W��z�k̤�ũH���F�#4�+��E<����+��G�&�u�"b
�g��r�Ւ�FG8Px�c�,:�����}��D���ceF��ӓՉ�OŸ �4�[��1[^��|4��C�O���<U6�"�f<��`�y��qᇕط��=;b���u8+Zǖ���j�� �k1��<N�=ZU�
��YL�)�Ilysվ^�k#r��3���ͬCq�O���� ׫� 
�Rf���\��X�Վ��s�{���u�[s���㮼Qqo�a~1��� 	u��צ�𮗨]�B�n\(�d~U���ǂ���d�\��xR�M��6�>`__v	�sRO�\jp��|�ھ��ׅ�5ị�]2bGG"�u{��@��η���ɔ�>�������L.{��ߎ[�<A!��#��W�~�v�� au�珠����U��p���]񊓱�}ny՟�����Wa�88��|E}s�ұ�9��sV�9e��_W���d"�L�Ďi׷�?�7��9����ӐI�� �۞�Th�,�Tr>��8ְ�K��I���z�-A"��� �:��Ҽ��>��_��<b�c�6i���yp���\�(zks�s஼ڄ� d�(�=?J�� �;�fT021�����}ӥ�xy�]����.jJ�ÿhWk�1�,�Y��l��c��>x�N�(-��浛q�Wŷ���J	���wSxm�3^�c�j� �]��c�!n�B���5���q���A�)�O8��#��S��dQ�6��_b���ߵ8[�p��A�����j���f��(_Xgɱ�κ�c3����< �El�V�<1���޾����X���v��?�Q,H͙5ذ9�[*QD�i'���L��s���*a�8�s)"TRk�ek?$��"���2����jz�=+E�����j�V���L�6vٯn���ԣ�y��͎zs���vM+�d�]�1F�k�ּ#=xu`��&M�"��܌_��e�=�]����Dq^iq�5�C%��|�q�^�q�c �<үQ�c5Z��J�[�&ïp���?i(���v��ٙ5�:���;���#jY�潽uM-F?��'s
�MGF�:���� ��J,�m3§��������4���>�$�Ky�ǟA�W�h��*,���G�f"�,n�:����Y�1���7_�L�߹���ƫ7��sn�4:����y�eԵo�t�C �}=�O	���5	��������1�����;������c��N��m���7Y�zq�z��ׅ�Kj��OlV����+v �J��m�^+X×D�U��k���l��Er��z��<��Gð��$n�����JGU��Fn�kV�M�j�l_g�*U4��6ݮq�.�7.�;p0��_7�^Kor�F�{�ѿ��-t3��8���K�5ӕ���SZ�$����w�$��uk�1�T�V�=̥~�Χ��w@i{(�5��-k���f#�������ۻ$zĚ&�A�]w�q>"��\�l��2�ƫ�@�I�z���ǨIm��ʀA�^s����yͱ�q��W��kgq���"�3�wĚǇt� �ݤe�z���3kDs��s�����G-ݜ�D�ʅ<צ���O���sec�=�V�xE&Y>�T�B���� ����:\��2���������M�CqF�31�:�Y���֯<��m,q\� +�z�WJ��I����+�
��6}z)�n~��97s�I�1������R��ߴA4� cvA���P��ߚ�����ݤ��O־C��>��k�������)��Ӛ��Zh�a cx�<+�Lۃ�w5sΌ�k������)
���^���ޏ�H�&uyZ1�K�ni��xoĖ�n��f�1?/Z��'�宛Ն<c�|�U{���=;T�:jT$�c��Q��\��?�F]�3�ג��#��muo��9�+6-1��̥���R��ɵ#�t?��w!]@�9��_>�bDj����� �&�}�+( ��5^'4�$Ջ�ƭ.�tҹ$g<פ|��q�4�%<x漭��:~�6�.蝇|ZIFG����h�e��G��˓���`���� c�?�5�G�GX�0�@��d�����S7�r�;��5ek#�� �[�2�۽<�Q� �0Ÿ���s��\��,�p�Z���ZF����8��tQ~�g]� �e���E:٢�d�� ��k�ok<e'?��7����L�-/au���ٟNٓ��?��?�P��7艒����x�5·��٣�G��J�)���C3{�qG��>�g�G�<�wI��E[� �}��.߷�qمy��% �Ah.� t�d�~��)?Ozӑ�$z� �� fOtMRN��Ԋ�5�h ���XݫL��'>��~<���;�ǰ�C�x��V�.㽎߾T����99-Jz��mRf#q�ӥ5d23��蕶�v��=�z���y%��`�Þk�����E�\��_�����ګ��`�R�b��3��	�>����:���i<iH����κ��Ե�ao-�{tBۙI��_=Y��]"�u�o�?�m��U�Be��*�W�+\��=���������9� �r����'o��Q�-�����|H�ր�Ia<���p,M��n�޷�k�IX���y���X����x��#� �E:�Y�`{ײ~�':19c���|L�?�QM<K*�(eWu�u�r��hǚVg�X�5�T�_���~��dq1��>�]t��w$��#/m�_�?a�|m�hWV�0����c�^y��f��k��y6��3�z����:I����5mFu��O��V8T�I��ϋ>�����w�hw6��u�ϸ�
�����s��|Z���v�<y܊���_+� �B<?s�{����ol
�c*=s�Z!��䐽�V����[��?dW_s��i�L��]G..����Tm��YD�>y9�����/�GX,� hf;q�Z�o����>� ������_�l�uK�s�,G��j�&�7�{O�Ҥ�r���^k���ƚ�X��z}��iI3 _Z�� �S㧆�i���q��M+#���}�͞"P����������}GW��{�y-�%%��5�x�C����"I^tS��z׾�kIk��Jƛ��{W��B�5+=��{�/�(}i��%F��j��V�_S�*IuZM���`9�5��xoǐ��;��.?Zg�"�96�v�A蛗q���3�:��ɭ]I�D���Uۍ/\��4�<o�̑]M����k34�z���$������|cm<���)�c��5TY�/}�Ip�[�%���	9�����;�ɯ��u��ۤ1����{|@����&�)� W�4�����V/cp�=�U �ҳ�ě���Q��^	����R[j<+ml�
�u��YX� g,�3,�yvl��|��o�N���6�w��<�жzl0i�;J��2�����\ᬹ^��5[�-vX��i79�;�5���_|E���g�Jm�>q��žL?!yH� 8�y�W�_~#Y7�m�Ty`��j�]=��SM��׃�Y�5(���m5N�KծX|���}?�y-�A��]���k�_xlݢ �3ӑY��e:/����>�h�$�{��[n>�N��u�i��.�Jt�6E��S�?Jѳ�S��O}�C���~���&r?cԮp���X��o��|�Rw,k����q|Mi����#�j�y��'^��:ܗGpܹ�O��*"�{+�WZO��'Ε��א1V<+��?��m#�V3]��p��G�=+���7����h�]�:���� �������Y��gq�.>eՓ�9h��(�|���S���N�+�j�#`�2嗎�5�����;�����ױ��.�qm�ʒ�`�<�ז|kK}5���19�u�M�F�ƢV3�*i[4C/��A `u�.�c�g�_���+x�By$�)�A�^��z��]l1��8�{���=C֚mvT�0*7B݉���"�J��2N���ş|O�� P6�Ť�p�Y
G�d��f��� �&id8UQ��z�����<)����ZX�M:�9B����G�k����_�H�K}OU��r|��㹯?�5�;v�?3|�
�B���n<��4ܲ])_3�qҼ�I�}q�?F�;�#���q�"�rh���?�����˾#v�h;
�V�<I��&]]��p��h�f�h�r����sD��[�~� ;t��W����O�]���S��_Ş� ���m�+�>S�}kϼi�f��v�rl~5�Ӳ��e�yؼ��z1?SJu	�����5�u�������\�2J�ea�t�v��Y�����gp+�V��</?����jx�z�V]�v��N�:� �?.�)n>R~�S>�'��I���h�.�}�ڢ��}����?;UN?� ]|��~�����W؟�n����k�	kɁ����3qsI�9��̀u���(�=i��C0Ƞ�Gm>������2Au ��z�ȸnW����h���'=�:�g���~f3��cI�hʍI��k]rTڱ�@�u��Z�`$��8y��zn��|,𝶽�1�@�.7n�plN��������D���֪O����kw��ǗX�
��f�$����x����e\�W��[7Z�Q��t$�+��?��@��j�,m�9�m�>����%YC�=(�ܕѭ� �h�pƊ26��� S�w��5�����Me���:��]K�z��[��锒�^��6��`K?:-w�flǏ˚KW�����;����D�ȧ�+���A:|�X�*�O�e匘��M��8���YO��� ��T�Z:v=��◇-Ԭ:|*�gpQ��0�e7����H��?ʼ�|�N�$H�}d���֟�+'�8v��wB@�*���F���_B����2?���N�烦�t�D>\��^y�;�v�5O+���� ���_������[��+�3�Vn�V����B�M���r�6-t��Ǉ<[��^�A��H���^q�H~�>!��C�����u� �Q��5�|5�ԛò�۴���ڪ���F5#ȏ,�-���3G�n<~5���kx�$�Y��;�k-���ֽ��Ks�~�$����>([���(�?+kK�[K5�Db�s�e|Y���e
6��Ҽ�Gc���w��?�bӢy����f���2mh-����i��4w���sZ���:K�9#�W�%�������b�2��`� U��7e��h���;x�+�����@���k�'�^������Z=�ZҊ����� �z��$��3�ט|te��I�?y��U�_�Lww�����::��	m�LE�]�G$t��G���C�4��潒���o}�_;�ʳ�k�� ��4�`#� y�^�>(;[*����d�=$��V��Tj^��K"���I���_
~���<iy!���1��-��O-Zr���x��O>�1}�$�m�I�¯��=൜�;o��.=����$z��v�-y��k�B��R��v?��í4����{s�ט��/��K����18�Z�/<L�˓&����� Z���R�n����CԌV�%�z�q	�3צ�G�xFi&�݁�Tv�*��]C�߻�� ��^��=mm�V|^�k�"�A�Ğ\��r����엚mΛe/�s��܊k
-ji�9a	���~���5�3j1�$��]�=ꔚLV�]�菚���ֺ,s����e��i1�Gȵ+��@	��sZ���G�$_�(Bs�x�X�t��n�7���8������$Y
����;�S5[u�BO�|���W�g��^/0��9�XZ���ڒ�x.O_z�6�h�{!p8����)hyN�o�60� N�����/�I(�W�����3��Km,>j�;H�ghmw�������G�Ws¾$D�xȅ�&2+�<�=��
,��W�|U�[?��vX� �w�נ�H�7�3*�����;��'C���ױI��u(�K������5�ޣ�F���G�Myǃ�'1�9#�y�Rតs�h�c�h#<�����_�.�%�A���۔q���%�R�e����[*�z��+��C�Q<m����sI�̛[s�B����@bps^C�hZf���z��s��GA�z����!� MShWq ��%��[^Iq9`r����4���S� �xT0��yֲ<-��Vc�9۟ҮZ]�xa��2�3��K�vwR�ȧk��1���C�PP �G�V�)lC�M��;s�+����{�M���@'?�_�+��}ff��s�x�^�-#cͫ����M{Ht&Uuy3��O��:�t9H������ح���L6��eL8?��U�>�$��~p����^j}�Έ�"��$���+�lh��v�Ȇ�␎��+�M��֮#<�����|O�!2#����lzw��w_�)k^,If�5	�:���_<�Ff��Pf�F���[Z�����us��s~����0��#$85�R���\�����B�ӥZ���h�n@�\f�.,�4V���PѨ�5��<Ef�QIc.[��]��6ǖ݊?<
�����������V�qR�`
��	�(���%���'hf=�k���<�෪���Ձݟҷm���ty���"8Ln^��$�o�W�|N�t~ ���p 7@ȿ9�?�p6�=3Z�c�{�?�y��>2?v�ö��E!s����Wo���O�}_��2��7�� ��q�wz�㴛�y2y�>����~���U����ɕ �����?�L���q�'¸]ҧ�ݼx�o�Xd���ߊ���ӱi�f=3m���X�\7��^�j����%����?�8u7��������]{í,�|�O<ⰼ���-Ϙ��q������_	�|aj�2���5>��6��o�XPHH��������į��\�d���'��#'��w�f��7M��5넶�r�n= �����<M(���ú�i,���zq�!/�3ڼ!�9���n597�˞��z�Z��5����Ϗ�Ҽ�Z�Ū��1���/�z��|�}�R��,8�e�Y��%vyW�|/u�ׂ`���]��=�x7:S�0��j�Q�g�6E����+����ԛ�i�i'˅pq��ݟ����|3oC�azu��~)��둾>P��� ������qw��~��H�����k���=�9�I���x�e��f��x�o�M�/e��\��� �����~�槩��yF����Œ1K��z3�K�|1�fO������-\^���/X����<�_Sx.TԴ8Z|��Ԛ[��+��Z�?�SJ���$S��s�U������j��X��y�U��,��Q��nk���:x���v3�NM��t�^��Y�m�i���{��S�;R�����L�<7��n+��|_L{��Due�X�� i�����-��gw��_����|0��<>���z~5�|HRтG���X��dP��^���?�yU�<������<�?'�� 
���[���'�J�2[���@.�#��k�#ԣ.v��3�7�Mͺj����k�5���Tq�_Λ�� =@�5�V7g]9r�|�o�O.5X��$�5��~%�-F�\����	��B�I�"�� ZI> �)�"p��Q����N�_��m�[(rIg�^k���?�$L��7s���+�o���S�r��_�P\��Ĉ�m� ��e4�AE��5� e�B�=E� �Gs�y��9qi&��I%G,q־�����'���Ĉ}\ֹ�xG��*�y�f�G�V��4������|qc��l�X�p*s㫆b��;�_FI��ˁ���Q� ª�`'(�w�����۟6��i�b����k�X_'�����S�}>�
���B=w�?J�k����%��v?1�����픷8߀zն�	��e� �v�<Qg�xn�2�=��k����ژ���gV�f��V`�r
WA�޷Gķ����HP��z��K�����1�����5��P��t۩(3\5���]L�t��'nJ�%=N�n��V淰6�pq����x��mA�#%>m�q_O��g±���2����B>�f9�Fz����a�a;G�+RD H��y�R�Z���fb};�W�'����%���c���_Y~���.��A��/b�{h�>l���u���  ��v����n�`U�#�ֽu~�;Tf�\G�*���Vm��� �:���!8�B�vXV���� =��N\`� ZϿ�v���;y����
[ڂ!2�}M� 	|$�%�Ɋt�n�E�fϝ�~d�����Fx��t�B%�픞UsҰ����Zn��&���@8�1[� �v���B��oB08�����v|��v�����m0��rP�⸋?\ٶߝF9�\����Yb�}�uc!��k�ּ�9����?�c��r��汫ʬ����d�t�.�J�W�]|i��A[eL�ɴ)j�4_���bF����N@5~�ៅ�a���}��G���xdˎ!�嫯ݭ��ڟ$1��M@�8��b��I� �+��K�ThX��i��_�+&���!�Who�,��Mbld�:�L��6�o2� v���}z�	�a�����b�'��O1G�*8<go5>��k���_�Sf���������~oj3��<�85�j�?HȐ�1�}�?�z?��m�g�c#=|��4mЗZ��w����G1��N{�������v��b8�W�� b�Z���Jۏ_,`
�f���χ�"�XQ#b�tG�F5'̏5��}sy��#�7��у_6_.�kx��h�y]������KF��[�Pێ�i����-z����0R�:���Of|����c�~1���P�l���t)�U�o����J���N��^�_�����x~ƿX���BڋEm6���A���\_�!��G.	fJ��|u��\7���ji�?�\y��z����*N"uԑ��qol�kw�lle���|� sy-�1�#ֽ�����_[�����Z�>�5�M4�>��KĖ�6+ߊ�'�.挡��Տ�Y��/�ֺ�0��s��� 7�A�^����fٿ��Kx�@y�CE/���?a���������f����~9�V�'�W����.	�_c�n�e���G5����u&8��O�#��r� �+�o�z"j�o1��t�|�y�9��{׀u,|8s?���l�m(��s�ֵG�=@���C��Z�+���~��Bs��7�Er~��s���M�����ק��T�|mᆒY#c�$�\���7���7�ܷ����b��oD��G�d��+�-|!���5�\,q±�־��]���C�5һ2��1ZTvB�<�G�� 		d<����Y�*�lv��<}�GK�.�s����^"���~(4�-�<�}�E�Q�3ld��o4D*��g�߈:Eƚ�M ��N�Z�g�� 
x�K�8����W4_�:�$��+�3��w�#��6�ujy7�h!�[i�P����Ew]�7 �Φ���Ś�-�F��*�~�HԼ���������|�q>.]C6�y�������  � S>2iw-x�kl���ʤ���[�v�gr8*�\5�9�B�NX��g⥺�EM�I�l�玵�1��_���x^�q�Z�$6 x�V���=wU�a[Y�c�P�^|��ΕU3W��b�5ѽ��R�n�P �}���O�t�[W�E^��k�k;�i�Qm�]��T�����K���� )�������T�h� ��C9��� ֹ?G�xOH����n�n�^����������Q��&�*~�p�A(MW()ug�~֒�����#�6w�y�t�Z�>��p[�U��A� �dx��M�e7�N~a����TGO�� X�Y���Ÿ�+��Mqz<����=��.����c�ir~^:ױ|-��hϨ��.��Ѧ�t8j�Ѻ<����1��u��N���d�'�n �ƹ��@�����;�%Xs�V�����Yٔ��r}��VG���k9nt�����Z��'l�	��s�>C\=s�� �S��X6ߗ��VF\��C� 	Ƥ��ٳ�4��#��A� z�ui����WW���x�k�MI[�����M_q���&���K�>TO;6�5���}iO��RÏ�"�$��Rd�x��[��w▃�nt��8������L>*�8"V�5��H��U��f��&�v��1V>��_�{��d��ý����5�F���BOM�׿�ql~�$BA�eQ+0���ۯ�?�e�h�A�qN����>�s� ]���� u���D���O�18��� .+�-S�	���/��W�z�����#��^t�1��c������{�����H��5F��� y-����������$ʨ��x����x/�"1���.q�iё��h��O�RI�mnsִ.�7i�k�ZF;��X����%��8c�#����z̨��kNx�#���k��]�l�f�z��~8i������rE|�������<����U��H��{����� W���|���ck�t���� �~��F��8�}+��-���=��f!T��׿'�q�� xrmb�&Y����Vr�싍'k��4_�vw�"��Ct*w7z]��uk��j�g��f�<'��t֑HZ|�5�և�Z.�g�����zV��]T�+9�|R����[T
���1YW?�m����p��d��1w���v��ƽ��?쭠������d���lI�XԭoSH���v����1��o^�!ү��r��ç�U����ţh���ʋ�m\b�I��6�},��8��A���:�[��ʻ^�8�\S�>?�b��+��o���Gm����uH�S�Z{x
T$z����Wdi���F���� !v*+Λ���p�T�-,����~��^��Y��Ċ2c
:����7_gݺH�O�y�����pON��~�~8x���� yd��g,D�
2n���h�[rI�K½E���4i� (x�Y��� �?C�M2�"��Ξ��y���^��M��$���&��cɱ�x��k3,L�;y=+��d���������{�ju�Ib���3�&�)�*������dq��ksT�2�D����3͕��l�i#���֏�Z��r�QZi�o�����I�֋3�Ο1&�����ړ�h�aG=i3�u� �y昅_z�<c�D��S�T����^Q� 	-��q�QN�l$������Ey�U�{T~}e���>�
��|]x�o��ٯ�>'���Z$�,ˁ�|Y�K;�/V�9�e`H�V8)ǖ�b�ޥfR0V�G�^Co�,����~ٷ�<�n�W�̏+�C�Ia!c�ڴ�ė�ۘ��Zώd�y�ޓhq��U������ŽǞ$%��]u[5U�wc��'��M���Q�3����q��v8�Z��+����C�5H})��Ԥ��h}��5&M�L�g�Ƶ��y��Z�i�k�cs���.�(�WC�܊��e𦄴֮~չ�<���������3��?�+
Ilr�6�2+��Y����S�8��G�|`�d�O:'р���S��m�$�����|��;�#��2����(7���h|V�<��e��@� 
�o�#C�C?��1_6]z�� �S��x�A�ʺ���>������0V����V�?<*�?�UI��_+[��"���R��ᱽ��EO�L�S�g���@�ܬ(;��*�>�R�s�#�W��,���?�����R���O^�{(��Q�c��:���
=x�_#��V��{��䖺��������/�<�6���*�Aɸ�Qh?4�;uY-VA��Ŀ�v�6�����m���+䋭H�+ޤr*Y��O��� x��WK��O�=Xk:����1a��f/QH��4g>��p�d���d7�ӎ��Yj��q�ɸ�8#ӥg-Ϊ+CV?�kSE F�Y��K�w�Vn�;�*���M���J�_«�
k%u�ZTe8�SΊ�5�ӷ֑�oZ���ubG�3֙����g�^���7�d�ߘ��d��?7�\��I�8��E��ݓG�D�^W6ʕ�8>�¼g?�b� hK���v ����o�G�E}^F�(d�@9�}�i�'ù/�a!K�y� =���6��2~�nk�+V�pe��Ȩ����7��~�i'��I/����0H?7$dg�}C�+����KX���C�䁁ھ*�_�(�A�ɱ���o��^7��RN1�5��׼{q�Hf��O�Vd7T$��׵?K�k}2�-ٖ1��9����3����Ď}��<+�]O�h%x�r�I�J)�sK�1���=����Z��LU������y�ڢ�\w�w�5�|�\��O�ҍ���00k��~�[�s$�>�9>�_��N���J���5Ţʀ�91򣈱���+�XUe�j�6��z`澗�ňl~���]�Iګ��� �k�jW-��C�ݻ�D����<.�t�l��z��rf5g��*��㷒V8�	ۯ� ^����6�x~��������|]i��I��ĸ⾉��7���P>����G�[s�~1ۈ<O�p��c��ȼ?�[��~��n��n�ۏ�v'�3�֗�um4�!��A�+���E^	I|Z��q�i�o�7�x��ll�����F`�[���<�\w�5�n�b�s��ol�uKs�E���vIʂ)�񹫽��ƙ��X�� f�� ����R~�W�G7���ڕ�r�Q�·ҕpm��s���oý"Kb~�_.��+��}k��{1�}�$qJ�\���h��B��W��Hj���/�uim��l���gV�E�e2c=5�L��n��M���V���dԲV;���-�X�bE,L|�79$���
��R5�yǿJ��%�R遉<d�*����>r'<go^kߢ�)��l��z�m�N�a�~���z�
�����H`�������]�<�1ۋu�='!x���=����ۊv��ʍ�c���1c�i�1�
l�1§'8��V�T��yVѴ�x
�j�ˍ9H��"���k�UI-�������Ox��G��o��U���nf���/$��@�sO�:����<��߅o<e�7x����&?�� �(����$Ӽ��[*�Rq�����9J��!AF6+^*�.�L�O��k�ޓ�3��}��?�zv��{�z#�X3۰R�9�p£��v�
[�!���F�fBc���W�x��y���{�P>�
��)�p�泵Kx�C�	5�T��9�c�[�z��!���Y��2���޾��7�� �d��w�u�$��2�h�V�)Os���1IU�'�V�<�U�.�G��Ѳ�ԊH.����JH�eM�bb�{���-��H]�����Ҷ��������Ι1�s���ɵ�I�I��r9� 8����@�PU~y��1�a��[���\h::7!<���c�>�,��޵ͫgbo�������c%�6�J�Ҽ?[+�ό�Mf���6�F$��u�\�nD�����V�B7�g��%��y�ݼ�=#8��]��/�.�|�u�����B� ��j�J��#�}��k�S��8��O���c ���H�ח^�,�zt��s3��� f{}J�]@ҐG@��6�t��BCx-_����m�-�ɡ�f��4��V���������T2�8ǭaN��"�N;/����i��D�&1�ܛD��lP��sZ�<?��� T;`���o�oQ�L��.��X$ ��=*牔�/��Gʖ����Me�fEp� t�� EO\W��c�*?�����grI��k�����u'�|S,B<F[���u�=�t�dx� �|'�ȩsu�Gfo���<�"KĄX�G��8�� �w�>��Z���c��_Tx_�ї�V&�Sy�ԇ�rǰ2�I6[��|I�߆:mΖ/-�V F~^��ۋ;�"M�U�9�_���������=T���X���ǥ~E���;-zp�+��w�p�ާ5h(���U��� M/jZ��Ih��K��.��QAr�����0>K����~���YE�w~ˈ���;�Iٞ��6�b���(�9�O�j������c�&h�wz/�]GĚ}�ʹ;� J� �� � eƷ��I�|�H� V�x� X��z��+SᏉ^��{�۹?�1���~�e|�d�eq��^��Lx%�;}$Dch�G�+�����kS*����������w���_��L0y�Y �_�5n�យ�Z���)
:쯫��f���m�Q�ɊB:�@�ֻ�g����|i�+9L���+�bfҧ����4�Hǰ"��u^���� Ǌ���k_�w���_M�x|z�	�S�R�(Dy,A����j7Fq�l�F�����M�Hx�N}���y�[�6K�lc�v�6��_q�?����Y$6��y�wa�=�X��� \|7�y���)��K2�2G�aC�����[�O����͂+�4p�fx&k��Qc�oH�a�Bֽ�����^	��|�
�~��G��-�Z~�&��I�!G?�u2x�f�ir�^I5���Q��4��s��� �cM��S������ͩMJW:�SC�<#�[=���E�v𞨳F�^�� q_#h��-f��`�Wq��6�#�Y̪:ak�t��:aQZ�ۚM�}�C78�kEo 8� ��_��^0�q�Ό?���w�x����G����G�%��[	2�k�u�F(n���|c5��<i�)X��@��+�����n�/o&[���*a�4;j��x�w�\��������5�3�GŚ���i(�8�� �_�7��p7��
6��]L�sZ߉D�F�|��{��#��M�n�A�5�z�_I�Û\��7#_K�>�|/�Z��0iv�R:�r��:�3�~9)�U��/9�xSV��GX�l�^��;�^����(}�޼~���Šo8/�{�c�6:i�QGI�Ch��[�SדR�Z��Q*�>�=+�o��9yF��g��5%��� B�GA���q�;F���z���@k��6FH�u�<Qe��z����x�MS+#D��a�)#���O.����gG�G���J�|���\��<Oe����㪰�9����+��莽�T�&�֥S��$��E��nz���^���R����׉�5&�&�9�8�b��W���%��ǿ��C��چ杅��g>ռ(��y�Mة�����*r��t� �F�G<����\��|H� �>��<ױ|)�[�{���1`�
�)�hr�i�C�>%D��N��� ����|L�5��a�k��#���z)�x�Ջ����Ź�M=x5f`)�R�d�zS��k�ni e#f⪛�.&򭑤c�U�xo�Z���ac����.>U�����ٶ����0��e<�5�[g�G̯#�<�?T�!���6�o����>�%��(��R�"�kE�}���|���Z�G;@?J�W�Gs٧J1FN��m60 z
��L�v���_����
�\����v�7�H��p�E>8]�4Puw����k��|�2�&�v��j��f�h�x޹��nIE�>��j��������=f^��qz׆���Z��yk؏�f��5�߄���ε�I��_^�*���4�I�o X���t�w��
�;<-����� ?+���m����Y�=����tg�V�kC��yw(��3x�v������ƞ�º��ce���c���@���
��%(�x�����,����W��+`�d^~��墽�n���kɥҼM�[5�Ä<1�����;�3�+�ְ6���k_ٛET%�	���k�~*|+��{�nw������~!x�T;-����Es~2�5�3:�Io��֎��7��@iz�����X��+�#��Isa�_+͊��g���:����߆�;�c�����x�[w�`W��^��R~���~�Z�͵�t��\��|}+������u��rO=ՎI/�]��<]<�c��9�ъ��Ɨ�Iv�W'�Z�I�{� ��㈼+�Ct���'1��?�}�y����A���� �����9��$������ȃǀG!���3�B�H<�;sJ�����}{��ڎ�����I��}+ᯏ_o<a�J�r�`�.1�z�C�O4�2�q�=k�<O���9�9ɭh\�v��x��|]w�O��[�#{�}kk�z��}�=Z`J�c���/�[���9��Y��O{un�@=y��'͡�g{�L~��� 0��16��p�{t�_jW�]^;JCHI��5�_#{�_��kǼ��s^�MC�ZE��.p5[p�is^�S�oݜ����z���oU|��+FUBz�*.᣾R���,V���a4��;��Ǘ�χmභKKpv��	#���^������v2�q�۔��Nq��zW�|}6��c����|Ih���e��n+�_1�_�������u�H"�I*85����&Ҽ3s�ʹs\<�u��^k��j��_H�7f���>2�' HG*�zZ�$�vDe��_�O�WzޛkX@ �0�S1�  ��cT���i��-�K�\�s^�_�����,�Sҳ>'�Rg�K6��k�Q}Ǒ~��4_�)�S�k����im�́���n+��e�Bf��'=��_�f�d.3gp+Ѩ�L���3�?�Y�?q�ؐҰ]�~�r1\'�Y�Oj����qö���F�ּcA��%�VF�p#8�y�/K�Hr�ٮ*7�H�Inx?�.M����6]��s^����eLs��s���L�d���t<\�ʾ�+�<Z�����?���Ǘ
9�� *�־5i���(RL�'��_2��IU�0*y���J�[��͜��DFZ�{է�[$!�]ݶ��_����\c�j��շ>1��ѕ^I"�����{��-|Ar���t33��8>�+���+��Wo�.��x����\�fAݚ���^)���A,R�ܥ�9�u�'J)�BRf���uU��&�U<��x�sV��uP�<�rſ���_:��N�-���N	������+\�����߂G����ght4jkV}�֚�nm���֝���Cj?�`wC ��q^����ڴ��&�z�� ��$�<W��׽��?�!� וn�՟B��kP�A� �U�"��Yc�_4x�"!� � /�_3��C[����2�q�9ϥ�5�*�I3���r��gf��U���[�w�31�3ZЮ�.[��q�
�F�ž1���hI���5|Pי�m<�����Q�4�h���+�=�7��#�J�%���[��O�7�� ��O�[i�k���"�rX��?����ůj[a�E`�p�1�zu�n)�8�Os�ִ���dh�Y�WpP�W��_g�o���>���?�Z����+�p�Ms� ����9��9�a�9�)E�r|d-�Q?.j���s�O~@�)\b�('�t�q�C/m#�#��v��L�~T��U?*�^JT~T֫�v'�3���4���i/�6]�j���W��)��二����wo.���Fkt{������
�Gh�F1K%���ӥ7ؘԔn��R�&	�U>���u��2[ld�"��߇u�Qi�tl��ld*�	�j�[�J�;KD2\��/�"����~��M&�M�˾Y���W&���G�����3��-�F��<
 b2�0�'�޽y���*�qV�R�0�  �⡑z�W��nn��"��!_�c���;�犙�jHm�2�3�T�Mkn����V�I݂zԺ}���k~=(�zz`(^h���B(�����F���^�FM��i`f�Ԃ�)P �눖N1Z��֡��qRI��zJI��Mp���U���W��ۮ��ֹ}b�:��,;�1yh���Ҫ��OB ��[�i�;+��6��Q�U�������5k9g�>|v󧅡:�D3�̭�X{��:����t ���玼4�,��o �9�gZ��k�[��Z&����	�2��矊���%�4Ȉ�9e�kCJ������⦺ox�O�&��[���CpMwr��-,x��]a4�Ua�y$k׼q�?�M4�h�"���汮>	�}mu;i���n{W�[�Vn���j���z�iT�QS]O��<*|7�Y�9�k�/��n�l��l�@��/�� iAw��}�8�j��u�I�*x�#�a^5{���i[��o~��������?����_|Dэ��#*�q�_x����ҵM�*�B�-��_|L�k�ĳBWk18�?t$���#��せ�-�z�7���m��.�&
Xey�񯈼3<vW�J�T�_t|��4��0[��]��&�{�裡���cO��s��S�@���%,��y�y�����Mi:����Ϊ���A==��O�'T�y�rqUć��c��G��6��w j���� �m��`����+��n�������Z)�`�����?����I��r��<����f�X�;����$���y�b�O���z߉�/�n�{��ߏk�0C� |��&�W�:��k��W��vQ|���׋�����ǡ�Ϸ�^��CT�4�T�a����bs�^�%̮xn:�O�||Qu����x��6��!H~R $z�I�X����	��V�����V���K���a��s��~	���?6'؝J��R��שi:|�m���9�k���~>�~����#�۞��>8��4�GA��2��1��W���s�g�,�Mi#���X�=���ܲ�F�r ��� ča|O���36fxm ��-�geTo�5����>��'�9�>0�#�{�3p�&s�կ�����=K�$�����]�?�A𯇭��bXu@�?�?�Ɖ�xR�6��@�nWr��緍,䳐��í^�H�Ph-m~idp��<g�l�R�lvd��Z�
/m�[\�;�Q����)7��_xO�n�&���IdL�˸��+�>4��|�����X��}o�ګ��W�m-�D�<�ӓ���?���֏�-=-��H>q�k*jQ�cv���:�<G��7����O�:>�S��\�O�Wr�޶~+xj�\׭��?4�)>��S���R��y�ֵ�@ex8�Xwڗ��@����g��|;��%ưYXd�O��)��.<�����ֲ�kC(�g��,��͎9'�gܤ 㡯�_G�}�A!�+o��)�~u��ī�1�I>���� ��ғ�4�ܲ됀����]�Ǚ�Y����y��[��*�I�v� ���|�R�ֳ��Ɣ��������Mo�Y�yt�<��*��^��Wh�����i���	P s_~���ׇ�a�Y��>�8�u?�*ϫ���O���;J�����jW6��n�A$d��x��K���^��l�����f�C��3��t�8�lNv�� p�4K(�hFL��I��X���Z�>�=�їWp�ӊ�,��N1�2��b����X8�S{�n�Sm������W/k��T�e���;Mz����$F��� �}�k5�\yj2��Dqz�N��8o�OR��ϊR����30�c�W���"�<���#2̽�_-k���Q �%� �z�~,x�}gMc+�m���S���U�3�㿉&e-!�n�T�o��{��Q4��ޕ�|�+�P�_{��P�+ex��(l&�GLW��<���o�=~�5i]m���U| �<?�[�2vq]Ǌ�2]iڴ�.ݪ��E��o�i������t.k�r�cĖ	���;lQ�wz/�j�+��[����Տx�Mӵ�.�峝�b�o|rx���� �\�S��>�E��nm��p�XL�̅Wо��H�@�Rw⼯�u�����<�ތRZY����[��H�T�tK��Af���6�ɒ@�T�򫲡i${�����˪�	�T��u����ǦX���s����c��m�� $��W���61�n��8���G�Q�,Q��Ȩ�����T�\T�Z��r��Z��8�����k��ۊe�����m�[��K�Ŵ�. =�J��)�Ƿ��R�r1LD�Z)��������^5��T"e�m�E"҉v� ��eȋ�3���-�����7/BhGq�PI�zޟ�68�;�S���W�j�H�?ʸgOH��=�z�3�X��R8�y_�?�*K��.H�z�ۖc���U�� j��F����.Y�
��Y�n���H����~\��>�u�܉"��;�����/� >Vc��\�;���u+��[G����=?�2xV�4��L���df�;X��/��Îk��b�������\ut�ޓ!��˧,���n��Z=z[U�m�����R"�:��^}���+ȓ��#�:�%�Е��S�Wː�;���d�s�p��<Wsߥ"�v�S�N}�N<M{j�"��WК��'p� f���a�0�u�^x���r�1+�&��I�m�N;����l��� yx�u,:M��Il�p)\
���� ø�R� �A:��m�c�JK�`��ϲE$a�� �O� 95Wf�ų��熯�j�%wr}+��q@���/�K���۞:�;�-�S��/��œ��p=1^B���?Z��^<�,;�E��~��ř���]���8�&z'��<�p_�5C\ԣk�l䓚��-��'� gҲu�|��g���R\ڝP\���D��XK*g�H�$�d�+1�z���k���r}��n߭s��k�qLG�pMO��F����JƱ���#=�T����Ƙ��,��Q�ʟ���Kq�{�������vk:($��������x�@�L�Ч%T�CShD����N=:	�&�ª��B̻��N3ނN�<U.�]�B���j�����_5�����_'�V��I�k6I���s�>��T136~��x��x�Ek'FrOּ��Oͪ!c������ڠ���y�6/=�9�F���>���O���1�l�Q����*� ���>|�@k��u��v�%�B�q�o�K��X6#V�Ep?J�8�� ��vn;���D���f˞�5���">�D0n9=k��ye��_H�v���{���w�N�ı��d*��9�+�?h_&�Pr�߃v&o[1;�+���,�&�p8����y���$�W�WRC�#��m�t��>$��{�z�� �L�G�6�|�:��Y���'����'�x���w=>c菅�#ڌ

�|T�f�'��� Z�~5��4�$ۏ~�3T�֟5��� �w5�V-t�s��_.b�O�&�e9�R����ɉ�`��B�"�F%�#Ǧ��Y�.����@�Q^���?�yY���x>���6��t������ͅ�\�&q�Wu(��5����̞&l�k��u�m�3y�m�9�|K��Ri�v W%�x�]J���#�#ֽ�Pj�<�;�t�nvx�UFN�Wҗ��f�/.y�����<On�K|��N<W�W��Pj�l\F$�n3�ק��*oc�O!���9��~�a�5�~&��x��K�9ё��n�n��q]'K7:����X��+�T��$���9�/����O}��Ձ*O���_o3��}z�yq�5�u�J���"����#s���"]+�V1,n���0?^�y&� ��R�Y�־|!��SKw�]��\m���+��/�[ͬK䲳d)�eOr��kҗ���H�񎴼�#�J�9����|���$4��<č�p���݀�}	�$�m�5c;�9��\��h3���[�o�^�w�~$�f95qT�o�RNb�^[�Gk!!V=��[(I^��t,ø��J����r�W�Ԏ=��-��go�1@))�_�MD��
 i]�h�3�g����y��❎A�ʍy�r*O,T� sQ9"��7~�N�|�խ��zT�"�K���q���v$�=뵺��R �ǽ!g�ژ�8J�5���+VS��ƙqn��?&[�y��.�9ٴo⼓[8潻��o��J���׉��S޾����>~���n?���?��_A�=뎹mў��u��a��sU4�d|Eo��PI5��y�{滿�����\,g?�y2Z��v5Z�ݡrϏLg隂��6��' �t;��IQ���-m�]:s�!�d�c���>S�M��E���|ض��01Xz}Ԗ����F�I%���:���RYD�n%�O$�ڵ�*�:����;]������Be� ��F�t�G�*[�Soj�`���!��=�:��L]��?�֯�p��s�k.Ue��s����ɶ�1�=*��OA�\��u `m�*��rA�Q�3n���?*��3��+�[�γ������ �Y^"� ��:�ג{֧�UVGf��������~]� :��Z#h����ko1W����V�������u�YM�#8`0Ҏ9�r���[�#n�hf�3�M������=�i�Z�� z��c�^Tr?��1���9����Y�j?ޭi���{A���qP_�<�a�~�R��Q��j��j�^�e�|�p:�M�`Ӛ`It�;A�����s���}����V�g�㨮fe�!����j��Û��V����x���rO�\[$[��ӏ�\�Ë:�?�zF�c�jђ8S���z#���y�xS�tߴKp˟�f��c6�}���ס�TեҬ�E�a�q\E��5;�%�ʳ(�⻡%c�qoS����I�-� ����7�����l�ֽ��ͫ5���`+���f#�,*���ֱ��8�­Y4�r9&��Ҿ�ף�ύt�Ἰ��ۃ���|s��Տ��*�gl�Nj� ��{��o�ɺ6$}������ϓpT�p?J�n�At���T'ޱ��/ѿ����a*1:�U����xA���]�����:|ѳ-�� �*�����G�5�o�^I���xx�G^Q:;��F��R����� QTG��_��랜f�uJ�F�5�j���p�KHMa�8�cE��/1�6�	���v��l7_��o��_̱DӶ�>n:�rc8��Y��Wq�D�#�l�щ��J�Ǹ��9��ć8��<��nZ�+𤬡��ڡA�ׂX���0N����� 	�ڰ+;o^��k ?@��uM5���#�o
�'����x��e?�NO�W�|V�t���/�}6����8ԤV�Zɞw���#f�kX�G4�6�{6����M�1����Rk+��zݡi���pEy<�/#�id���9b��&���\-�/��5���y�۪w�W����`�*��h��|t��-�!�z^Y�_K�]4ҝ��5ޙ$�sҝ��\�D�����QP��n3���:;��rޜf����r���9�U��쇧�1����I˽v�W�?������f��\������v@5ϥTh��չ�	��X�7WΞ�gY:f�m��ek�~�z؆��Rž�9�g����j AV�_���zS�6�5�^I�ͷ���E�ݞ�� lS��ГҐHs�~5$ ��Q�n�R�Ȥ'Ҁ � �z�<um�$�y;�U� �dޯ�޶&!���Yz����#V�ff��\��텎3��]���~��r:��6�q�:�/y��|q�@��A699��ۂ{ר|q���������y�dF+��ݤ|�W�ȣː�WQ��sNp8�\����=1Z��
i7,��~S�+�����Ĩ���w���^f�[����&MZC!f�ֹ&���02�t���"Z3Ԏ��o%��ێ���R	7�Ʃl�I�L��<
�?)^�6[2`�{gҪ�A���3Y�6�P�Z���qy�z�Z�g�}���-�(ʆ�{�~\K�U��^�t�k$M�gQؒq\�q�3~�d�贝B�HX�gu�p#�+� �r*� ���`s�S��o`���2�c��o%�.�v���5dO�=G�V+���sּ�ݳ�+�׼Z��b%m�`���s1���6�+�q9�T��� Ll�7)4=K����?Z�PԾ�3yc��oZ�f��o�ˑ���+Q�B��<�w���f}s��jU.r�z��؇Vkx�q���:2��cy�i2'�ң&����
b5�Thy^W�Fڑiy��'�z�CH#�$0>����cˌ"�Y�����α��5�u�)�����g� ;+���2���\���t&�ڴ�D(����q�1����?�y]R.�?ʽĞ �O֭���5�:�Ώ2�;���kU�EΩr%c����z4�̎:���"��6� ���(N��Q]Ǉ��X��J��eb;���wE���iP�IYTz*��ax&[�\�I'5�#9�3�.>���׆��+#��|p��ב�����KX�$�?���$��\fL�<�k�1��ɮ}��9��[�2})��$U#�X�m�*݁ɮ��9�u�6l����X�P�3�T��|N�{�e��a^��=Y�p �W�j+-�]��T����W�S�r��0����Ů�yw�%�p��	�t�A���<�DI���[��}+�BM?����׶xO�3�I v!O���g7C�?��:��mR[�(�o,�
�|?�]j�0 =�޾8]B�<��H?�?Ƽ��̞e�mioN��VӘ�c�*6�O��!ףy"kxaQ���G�y���3}�������j�9�_[hwMo��q�W���Ɨ��x�Wf��S��Ͻ(��C�MV?�F��227|T��m �c"B��ν��%�p�[8��;Տ�Z|Qh;�`���� 
��nVF������͎�pkY۬�68\�k!��(�z��j5�S��k/zǵx�^�!�]����u?����I�2
�/�~�|U����;X��'s��{/��I�k�����YI�ť�,<�K�<��9N��l� J�����GѴ�qa
ƄpV����Ʀu��J\� G�:��c�����ϒ��kH�2d���/����-������;�h�����ǜׇ��dvc�Z���ּI�$�3Eh����T�M\�kῂ�kQ<��0�n9�q\ޟ��6K���®~\�#���~�Ӽ9)fڿ6��_=i7Z���p�$.���`�WW5�G��T�~���k-��k�~^8�O��o�?6��{{W�x���|#���9뚛�`�0��S2>��V�p+*���BVg�L�`��B�3�>��ݢL���>�"F�A����z�е��֤i�1�Tl����y�{V�L��CRP*�ԑ�ȩUU���U�R�f��_�+(�
��0#�E+6�(��ҍ�ML�OzV�q�*
+=�ic��5:�#)�1��$��?�"�¯�' �PL�W� �1���o��ޕ���u����p������>�����<�_RMz��ars_8�z�p��&�_�|��ه����ZJ1>Y�ޤ/���>���O�'����#��q���rI�MQb7��<��#��.i�1x��X����B�2���x���ǥrN��:hȳ�{T��"2/�����VԾ�1���a������<����3�{�|Q�k��W��?Ƽ:�������ؔ��������vf��MǸ��<7��pӮ�.d'�Wl*�\W�wE��i.b�KvQ��.gy�r�O	h����3���'�<�<��4߳�{��ݫ�a�1���l�9�7�W������l�*W�(xyZ����C��܌���,i䡕T)�k����fI�M{V�l���_&=9�)顼{�����ie��� wmB1��-g݅d
q����/�����-���n�J������T�"�܃]t�z��u��UY#fnGzض��rݪ_�.�OҽE��U�Ny���t�Y�t;󎵻=����WIӼ�Q@��8�J�\w:iTS:�-$�Fٖ۞��jwҖ{v[3��3]��cv��wqɮ�M���ՁEbGJ󯭎�]��Ac%�� �d w���׸|F�`��ic@�r[쑆���Щ�]&TV`x<��	�=�n3�U��~���k��o-�hʯ#���ʬby�����D�b��3$Է�V�O���9;Ev����I&��3�Q(8+���ObŮ���
o�n ���󫋤����UN���k���^\F�x-�x�����7�!Ѣ�J�kv�Nfm�ǌw�cyX�KC�Z��*�1���KHٸ��{Ŗ�o��|�<��i#���^�8�}ir����c+�'�*�?2��*������������ڻ,�:SRD��v���OPA�=��~j����"��§~a�k|�;���~�UA$�~���V��2[^$�2��K�/��_�u�����O2FN�#�Cӽ}C�� ������˻R���H�����}��r�Z�a��\ O�k�~9~�WZ��q�C!�O��  �8����Sލ�Q���[�<a,J���0�־��g�=x�Ś]���h�2N0���_.�,[���x���/���e�����8� �[ c�i֕�q�V��?����/k~
<@�����6�+�ϭx�;Ti�ݴg�Z�/ڇǚ��<A0��`.v��}��#�'��H˖���Z�{2,Դ>��~����L���
ǒFk�OG$>$�d��O�� 믳|�{P�<(ciU�iڠ}�Z�������~�<������r�m;ݟ`�����+E����{���+��/�?Z������m��,B��3���<��W�~˿����1���yڌF>U��_��K�k1�y�q�
������k
k�ܹ�|GV�\��q5�gn..#VL�+;n����� �\�p��_��}%;(�?[�>���m7��L0�ƂA�� 9�����!��)����S��uOM7�����r}�գ�C�d�NP��~{ԸslO=�>�����-w�� �)$���%Yk��Ȯ�p�?�m������nLqw�X��Ù�>�q!�n�8F�R�.dqVQ-��~i�e�ߝ{Ǉ~%i��b�Ԩe.���xD�L�'�c��צC��R����#�+�ZK���omZѾ.i�(�ɾu+���nǯx;ESq,��Fs�_#��u�^2���py=���m�׋uA�; ^�����Ӝ�*|L�[�x-0�;sҸo���h� ��|�x?��o|5�@rI�.��[�m�Foү�J<�q�,�g�¿&��ڿ����>`8��_#�Ϳ������YG9=��='P��%n�|�j|�h���ٵ%������T`�1+Ҵmǭq���+Ҭ»���¥O�r)�.ϖ�L�o�O�#�1�ץ V�Xq�d S��P|��*�pjM�lzx=* #nA�����g�8 �E V�l�Y���̸lw���J�@���XZ�Ћv[�V�����y���U�Tlc)J�9�%�J���ɯ��5��kZ������e���,,�A ��E|��޾�u$��'"��.fy8����7sQ0�f�cw0����E����3Y� ��sҴ�z͝�#�֞毅e�.��K�ƽX��b90 ���-�n7(�	Ȯ�a.�Q�k��S|�=�<�mN�C���v����<i�,�+d�d9�\�ԣ�PCt���x�^[�q��qXQ���՜9t8�����`Hӹf$��ৌ
�6�j���MX٤��p=���Z����'psK�]��e���0
��j���0	��MQ�ԑl��$u�x�+i8>ƼJ��)6z��E$zf�6�V�T0�{�W�x�n�$$ Y�Z���ס5�j��_�oc��k�NI�sb$��'EC�4:�i�(ix^��{(�X�Cw�J�H���N�;Ԫ�+)�hn�Fps���Z<ѱ׆��{W����y�:�R��#��H�Q"������V���Vy݅���	ҕ�=�V6�g[�,%��[�ח�v���KIӓ]o�5�qa��H���w1�{W�F-GSϫ%'��X��nhT �i�9ԛ��ա���$gf�OZ�hňX��qڸ���j��ᱍ�y�LE7(�oI����$�����Üps]��qn�)�U�y~.tRwrjU�,A�ύ9�{��x�P����#?�CO�I�^^5�ɑ�w�k��8���.獈wZw��}h�-u����m�{�Vj�� ��dkO�?e&�mݎ}�����>�jbv�s�K�%���+GԵ�Y-�V%���B�$������Y�nW�S�v
O���x��D��� "R�ќ��O��v����:���'��� J�Z�-X�X/ݟ�P�m�yQ��/9���/���X��7:���a�e�@����h/4� �M�H����'�jjk����$;�9�����B�w�Fx2˘��a��>s^Y�E�׼I�l�̄�/�5�?����+��!^���?��|EV��
q���2^�Bm�gk�	-��>�O�@�2p����5�ϋ-F���o�`$+�z�_]ϥ���v>L�-�ϵ|u�G���%�S�,�ϥe���f�Gѿ�����n�c�������O��𞕦۬�j|�`����_�˫���f��8 ��Ҥ����bK�(�|�j)�ފK�>u���Fy�\V������1X�>ˀ��{VΑ$q�D�p��_Y�C�+|g��ک��r����^���7���u�\y��c���{��5���(�E��`s�v���x.�I乍��v��}1G3��g���{�hF��A�P5�.���H�b����?�@�7���P�Q��r5�=+Ikf���.�ֈ����C�l�[�hH�5}i��z���ћ�����t�j*烻#�rԵ�kF�L�`^@=8�k�����ݷ�-���P'�My�yw��j8���l��צx�#��g5�� ��x��=Rg�#����ݭv+�����K�c���ׁ]*���ɯm���,tִ�Ԣ����0�+{涧�1����w��:�[�U$s־��w�H�->��L�\�k�b9LlNy�{�+�Y�<�I���	=+�EIs#�W����Qܠ*Et1~�J����&X�IA�^���n+���J���e���R�,9�#��O��X�C|��zT�w�2ܑ�1���>�U��u��#��⓮EJ���
z�9��(�5���> Z&���2�H�z1沮<a�٫n�1�4�O1y�b{V>��Cg.��k����Ym߭yα���=��m���1�R���	Cns�A��玡��i%]���4�9��o)IK�3��\��n5۩�J�2Mz8|3��8jֲ���׋e��'Ϻ>���3ެi��w^J�M{����M�������b���5dy6u��/���TY `3��LW�q��ztӅ7�(�*����i��wGY�o#H��S�4�g�g]H<܃������m��{ ��*���o��Ϲ�H~囟Υ��4�9]�|��
%���8e>ۀ���j������0�$��|+����� J�k�4��5Iq�6]��ֱ�eݐA���~��L�_��lJ�s�8�=p�� �s��E��
Z6|��/,p=�Hn��#8w���c���b�q�~a������Dd��3��(����>QW����?�Z��k���
��٫�rX��Ē�����Ƶ?��� y����zP��1��Lx'��q�m���~G8����77��@W�^"񅿅t;W[t�����k������j����G*��2{#�?�X���t���� �L>x�8Ĳi��C�ש���]��k����s�֏�.��o��G=Ԗ���=R���G�C���x� �t��z�*�|5��̓��W��ƛ��fm>M��!�u��o�I�3
+�j��3����Rүt��mq$���z�g��z�b���gC�`�ʽ╤��uX�#�� >��2����~�����/�Q�z�.b�Y�,�Y3��ɟ��W!�=�U
�27��z�~���Q ���'��Oo�D\8�Œ2&����Vg�7��j����`��PI��ѩ-dPvʐ?:�H�2k��>�p��6~x�w��g�O�l�3�F� �dR^��I��I�/��!]���@@�[��s`�r�����$ y���︓���^��$� ��W��\���� g�I� ,�^)%��|Y++��b�U� i	���u�R���1h��� =��T���G���>.*qj�����o�(?�{����#�ҽb�A��a����SO�R99dP?���g늗ʴ����G���	�;�i�$w�b�^����my�Nw�z�S���x�Q|b1�K�v�<a�Mr,��$������|���:���R�ʿĽ�+�]�r�j�nZGa���n�gY���H��?���2�Gʫp�Uk�Ց�#�}k'�_	}���́x��s�������!�Z\�.�l�WMemá��p�� ���ZiP�jKŌ�p:�J���Ӓ����c��m4�� +Ҿ��4��7�$�&�~������=������ߛ�����v��#S��FaUwO�|�d�V��CH#⿊��'�6y��s_l��:]�ǃ�ٛ-���W�2� H�D�#���[>��O���hl|)op�T?6?u��C�-��N�g�a ��Np0s_/~�:]��6���,^n�1�5�?�'���=68��W%�<�ּ������;N�2���K�v.~�Y�m������X������lZ�362\��+�[�i���=�l�^zW�?<S<�Ȳ�r�A���~U4cf-mz��t���I��n	�o��w�� ����0v^�W�~Ϻ�����s2�`s��?�u<E�^xvT��X���ҍ�A;4|{�:.��Y�g"���*�Z̸�e�gC��$�ƴmY6|ǩ���SK"����|?�|I�I�K%!N����q?��b��w�v�n|�-��wX�	��:W�� �:���O23*��f���`˟����2�q�3Xڟ���2,�"� �L�(�%x��=���T��X��~,�#%�â��q�&���R���$���"���6�֣|&�d��d�Q����o�It�E��M#d�	�S������y�[i���T*A��)�E-���Г�/�-a[0�i�k�����.���z�c�~��T�)㈵-���?6[ס5�|q��֞ߺC_�^B�n�\�G�j�	uMJlh)>����6� �ר��s�����b�`��$�>�?�h��<P�[����=���'�I�-���B<�\���&�|��m�ښ�7]��� Q\�k�,��Ccty�S�sϥ_�Y�曧-�Α�Ej��<{���K��1q�8��^	��·X]ެ��6Z�o���hd�������ψ ���� wW�x{������U@���\���bvR�������;|ӟ_Z�t�^��U��־W�Ϗ�5{x�)����Xx��<��ּ�nwFI�B��2��E��:W��?%��#�@�t��P�hǘ9���/��(E�����V�4o����f��Kl���W����k��[1V'��x��^E��[E|������]L>V�J)�B��Z���5��<�ۏV<��%�L�d���w^;{��L����� �^}�?��O0BYm��vƄ�s:�>��5�>7i�Q���xǎ�4Gk�Z�#��x��>+_�@�H���=욄�һ1��ztpj:����;�'�޻p�{'ֹݹ��I�����ZCp���^��VG�)JZ������ʱaҽ{���曡��#|�Ͽ�^���8��g�,&@�<��J��ꢮ�q�?�|a�i��Ҭ�/e��Ƒ.I�m� xr�l���*�BM�l}+���#ƚ6��[��i_\6�x���dt�>��ߵ����.����I$d���7q�}+ɖ&Q�������Z��]�+H�VBǝ��#��b��C�g�[l�Mr��bEzV�ws�ؿ��0G��p�"���x�R�]*K�� lL�ƪ8�fK�ٞu'�5�m�Y=�qO��:�����<}�+KP�լfQs��Y��*�]�l|E~/E�ɤ�<���J���H�,ѳ��-źM���t�I?�z�6��{��G���X7Z�c��>��;�)�n�2We��̀���㍆�B�%LKEƅ�+��x�O�Ki"��	 G	-�=�+�־�Z�߄ź�����c�i��?�����E�h����ح�p�$Q���O����<1m����Q��d��2�e�# R�yɫJ�b~e������y�P8L�>"[��4�P�NCg�|!��P���ŤB(1
: I��-����劑�נ�S�j����E�U$��
�e��F����U�[�D�� �/�Ҭ�~m��+ؿc���Z���,l��}r��ѝTR�=z�7���tM*3�}�sZ_e[_�^.�"���M��_/�8��|F���Qu�e<�ާ�{�E\h���ݴ$�����+���s�<����O�?����4kDx�;�u�A����A��� ċ�{g[��!�=z
�{����5/xW�v�J�d8S���|)���^�Ĳ��f|�z8X�����\��ջx����ό3�;�Z�ڻ1Ӛ��&�d񥢠@�A�pG�kC�U��E����e8��]�hn�}��� g���ދ��f�<C�Mw?v�C�s_>�kᯍW[Э���f�mO(����\'���&��1��L@�<�gֻ/��k�+�#���^%Y���z��z�~"Yj����-�c1�x<�"{1������/�򡁗?����Z�/�o
�!T��ڼ��O\�ޣ=�����v��E*���N60[A�w-��8�g�R���8� O ����W��������ay��<��1��b���eo�D.�B��j� �^��H��(f���Z�6V�9$=K�j���m5;O>���~lu����?��� `��@�_5�~t��#
˷��VW���a� �/���ߊ�*�?�}�M��s�(=:�_r��_�������Ӵ�;N��K�q��bX����x��Ú���v�������|v���x��Z>�׌�ܣs�����UC�i��2j-hywë;-?���w�y���g���<kF���cr��\w��ψ�9�g=k�>'xn�Q��'��dW<��"��շ3�[���$^"�J�"@�+��%�[_Լ?�K�eg#�ײ�S�.���8�m�U@�-T����d�n�i#@��ӽ��'#�G�W�ԍ���)_�Ǌ�?h8Dz���+��_�	���R���W+�
�O��%!ծ]NW<j�+ꋧ%�p:|���SҮyM+�/Q�g�4�=��qO�.��w$g���*7}OA$�64=F�A��H')��Nk����{}h�f%�p	&���	�H���k�,�j�pM��RiXӸ��I��8�<�]_�|Y���<Ir�3��k��Еr�ri� ڮ��)�}]�w����~4�N=NkO�[㜧|��y��ls��4ּ��1�qBK`����ǚ�B#y��q���� k�睥��沾�͖ɩm��������Q�tz�q���;�R��*���]kd�%�Nk���/ma�7=N�rJ�5	����E^��7ínI��s��m�<+�bG�K�#}���V�gg��o͌��9綧�|��4���,���s7�����ӭq'�p���1݉�WU�m[�2S��1���.>�༌l�&����]�W�G56��ү��~�>��=��� 4�ā#0��k���g�v��Zۢ��01���s�k��I�������x�dQ���y<qa-���PI��g�Q�g���� f� ���� �-������W�;U�B�E=�{��_�Ro�.�^��Cң��|��$1�189&�+�I���y�/����zW���S��Mx$�<�^zW^��s
�H���t�x��f+�bMǅ��k���N
�� �5�~��c&���(x���V�жC�s�½E{�y�)�� ����9�L�'��q�l����s���^��B|*�o��S�3K���(��|��;�_���^{$����
�_|F��W��y"�׃Z�w=Hr�z����<Qk����*CȬF�k��2��?n��������cL.?���f��	t�Cw�����u�����ycc�m|�?Lӣi;�����D��/.!@����Gۓ���+��1nfS���?�q��c�Y27��O�va��<c�}5=���|�m>���8�3�C��|z;�$w����5G��8���}�W �y�S�G)�Ə�#IգR�(v���<�Mk�YMe� � z�=�|Q�i�6LY:�[��4����|�����:X'}���F�ⴲ�x�PWA��O�~(��߄�fV��ǯW��N�t+E��I�D�	�O��7�'�ھ��ԧp��N澹���f�w���O��W��*ljs��r~�� ����q����S�b�5(��F�t
I�k��5/iX��O�9d�PEy���-���v]�O��X�@5�^2g�5�I��y���-s�~�5��6aRM�/��7c����i3xP{y��W�|2�ѹtfQ��VO�mlm|P�\�g��#Ҕe��q]L����[%��H#�v� ԟ>��P�m�sȯc�/�M.ⷂ0���8��C�����.�m#$� *�N\�Jǋx9��fO!�5�_�|��J����|��^&~�^��+�ۄld��ª��Q��{�G�$��RB���/Z���q�0��\��+��[�k��'�v�^��UAɯ����=�ٞ���S�?��μ�B��H�QV��>7J�<���3>���~�ա��2����*z�����?Z�S����7.@��	�?�z�������%X�!�8�qVz|�"�p�ȢB܅<� ]���:ݍ�V�e���� 9�Zٙ���\�}������~��ԣ�����$i�tu�0�F�.����\i�`�c�o9滽
���"U z��X�:!���j�F�3�{}j��/�'���)h��U��`6���Nq��Px�T���e
v�'Z�wRV1��_��r.�+��۷5��� Uf�P��)�� �s��js�}k_���[b3�e�Ӛ��sʞ�>9\��M�a���+��k�����gfPWo��]�D���鰎~�j���$�9�Y�y=k�'�ׇE;�z��EpH9���`����V�B�;�x���6�L�7,. ���9�;/$��I��  On���H�P>0�w�5t��vt9����O�O� 	$cim����i;�[QZE�* ������O|��'�Tdd��{Y�GS��lu�:��o$�?� ����I��푛���z��[�Z�� ���A�_��p�^���G�һ��j�3�M��!p��$���V�i�W�޼CI֎���G=+����&B���V����I��� ��s�2`�Q޼��l[U��ۂ����Wc�쭼7�0VT*�=My��<mcc�K��*��� �Ʋ�i&�U���Z�wP�!I�'"��%Է�{U�##��N��o�S�vv�"���0���9�����j�_iUE��c ���˥�{��=��\\^��zd�޽7�7	o�2��� ~U����^���m�cG�C�2sV<)����K"�>��8���vEk��8����#Fq��׼>u�baq���\ψ<A��+����V����P� )�qڶ�O��c9ht?����b��Ў��<-ž� ���2}�I��w�}A�*� e�䯠���^��<Em4�U^���?��^�Y�K�g��/�k��r���|�Hح�?�F���9�48�|��$�i�|H���+p����o~#�	>�H���Gq�S���!� �����7�
>`�X�n��Z�SG+����k��	��O�qi!22e��<t漯�&������#^h�����GsʹV1j
3���Ҫk���w�9�Ԛk�x�_Z.��<W�[sզR�C���u^x�F1�������5͉s�]���3Q�nC���j�:l�1�T9���$m̸�^}�ZO��ӥIok,�Gڅ��k����mm��`�d��C`ry`�9�ֵ�=r��(���$�Zm��]������y���9E`T���p;M[\�6x@�xr��\�,�Ɏy�1��I#8��Gp�f��On�z�89�&���0q��eD�x�<֛"5������kzw��Ue�Au;��"��������������v��,dV�W�k�~"\_J�|�e&��O�=��?�nn�w�����
��L�LP]c��+���D�o��Ӭ[b�p�z#Y�������o�~U�8ɻ���� �$�!�8 ׇ�V��������s��9�}/ĳ7ɯ���sҼo�梚Ǖw*�4o������9����=���n4��yjq��=x�+���լ��.����g�����bOM���X�\3.��n�}}�ҍ�8:���X����2;���,t���<�|{��\��,6�D���z�{�Mk�����>:�j��LV=�<?i>A9��ٮ[��ll4��<�n?��k�����?���� � �`�Fյ[DRjR\D� X����Ӄ�.F�T��X�q��t�dq��u5�~�k�F����~s^��X2���� �~5��{-s�##���'��_֫���EvyuoNӸ��=kCO֚�硬%��R�pE�迷g��c���Eb��yW�G\�W,֧�JO����8��G�s���ߋ��L�=�����$I� ������w��f��Wc�v�`�m@��)�3^�?���J�j�۟�ׇ�'խ���8�_��if���`��޻�އZ�{�ދ��7�Ӷ�
�	��s_'�����Z��wV?xױ�o⥽Ƒ����1�Z�� [��ƺd�O!����T��
��^�w���~686��y�G�|-�׃�� �fSpY��� J�ui��j'�9009�r|�.��e�؋q��z�ī�D�����Q�\v��h�w��2���'޽�O��)��}"��$����N�*���#�r5R����Eh��0��ӆ$u��9~�7�;�n���g�Ui��?��G�c��b�\����U9O5������ )�`����:��Yb�Ewa[򯡿�V��y��9
I"�����K���8�U���Ɗ�֧�j_5ˋ_�H�E�=y���HR������C�{��Y��x#u!����� �@0�!=ۓ���a̷>~־(^�OM�i��$�^��|X��GHX����?�?CZ���¬����i�{  �^Ǜq�k-��d�M#��3�y�k��J6�^��>��&��_������ќ�uj���d����Tf?���K�cks�>��j�q<�g����t~<`|Sndc��kټ'�x�l� b��p8)���1���p�J�n�z�N�=u9����� ��\� ��a�;	��>*]B�lk"mm�{���K��<J�1�j�]��H|A�B�+�6x5b?�p���5L�H�Ԫ�� s_5��\�=�ly� �m^k�3�$.95��7��!����>'*��v�+��jȺ���⾛'(�x��gc��m��׭n�5����z��|3h�l;�̠מ�N���1^S�������?M�#�|�`0���+��vڜ<�|k$�yPOB��_���6Ny�m{<?��롼������%��muUO�@y�C��P����M�Ʒ6�v� 	<�����Q�Y-Y��IRk�Wㆻ#~�B>a�B�R^|f�g���
Fb��p1�Y}^�ԑ��|��-�w� :�?�� ���J��+�����%[�������R� ���l�vh��^���Tm�^�G�����+s�� ���W�-�	����ש��?1`�$��yG4�^4e%4��%S s�P致�����3�do!Y�����ZV������Ȏ&8�`g�y��+��'�ѷc�<���5k��������O��7ӮkE	ɽ�����oG֖�Rd�i���c��Ů��Kx$u�S�}�^N�� I&?��|p|�W�����ƴ��y�έ߃ZF:�s�[Sܼq�n_�����nR\3�<t�SxZ�O��4wK$����&�>3��P��V#5�^|X�cԌ�|��?έ�W�=����%Ρyq�#8���׏�p�"�ק�r�o���Ց��q���:ֵG�/$�G%���[���� H\���w>q�j��j��䈗�/�U�4&m������G}7��20A���z{C�����z��[x�:v��i���)���uV��_���@q��})�kv�KGx^�U������8��*�I>F��>K�[�Uw�<�Asy�����FkM,AS�@O kb��C
���4�ֲ�$�����o�/㸘�iU�"ѣ�I'���"�� 8��.1�H�-��ڙ��y�a�w�:U�*�,�kf��T���\�&�4���3�x�M��z	L�8��tQ�«�:߃����:���6{5�p�{Wm�Ru�A�J�O��I&� ����=�h]�_�w1X�$���a��ײ��>��4���� �c�𿆺g���mѣ2ȍ�eE}_���ε�v�9����l�G)�3�:(y�qwpz���o\�w�3ӥ}!6��lr4�VfBC)W�^<��קf����m�Zޏš��=��y�Y��.q�g�{V_�b�2C�p0H5��9��k62����D.�v,~j��su>v��Eաi07;�+�5�<G��h�.dS��>��*�(Ű�W���>�Vh|5m#�q�������z�Lv0m|3��6�O-���;}k�ε���-im<q�ڦD���S^��[H����t�:W��w�T�����T���z#�w<�἞n�����J�ߋ���Ð�_f���@K�����	\G��^�癈<q�x�?q���w�Wa�=��i�w`��j|+���2Kn#�B~�O��L�?i� �(�I�N�V�>���Et;��m8���a���<n���z���q���W��0!u���ۘ�θp�Ţ��t�n�	�PH�!,͓Q������u:?¿kP$�Z�����#�z�H��\��4ڤ���+���19�tz��]A���o����)����I=��Hݷ���%u#ޝq�{�p�G^�c�|A�kjD���kGR�7�iq��I���&���Z�`豍[X�N����_EB����|����۟J��H���֣�H�-��9�5��2Y�k��P*ʣF����i�<�U�$}��8%���x�eͮ�������O�]���/}w&ޞZ��9�'�_�v��2$���6O����;N����<|��;�j����lN,������^��O���!a'��H�sS�o���Ԋ��S#�ɞ��oϢ���֟'�2�m9]q�`� �疙��n ��ndfPb$gp�R�;��䏠!���0�����kK�G��� Y�.z��W��j���Y��U�;{����E�N�*�;�T�k�ܣ���+l��W�(qJ��+'��& @@��:6�Z�o�H��l�r텦6 ���v��aO	xw�����r��������#������J�95vfx�^��v�+��?�o��ӗ�Ksh�l�z���:���ֱk��%1��@#�]��=.[b�B��s��G]���K�F��m�P)=�
������\#J=���Jخ�jѾ��	�~�k�*<�\j~~=k�Ǧ�dz87��G8��xS��_�(��Z�-?��ѫ-䍞H��~i����>2W��ƾaҗD{����M����&b�7�
>��	����L����z��	��J�N\8��yǯ�^A�-�bz�_S��P��r�����^^Z���b5�6���G�0�[F�q�}���mj� l�����]O�-�?mG�`��9�ֽ�y��\� ����f��(P��;}j��>�y�SL��O_�S~��+��e�֢[ɘ�L܅��+��?xF��4�@�����yb"��cIRv��t��L�tq��A���c��6�0:th�ᛟ��y���q!��A�Տx���ձ�_�\�AƔ��o��\��X���ɨ��}Z����� c�z\��U�� {��3ȸ%�h��2���r����o��AVG���r-c v�xΛo�Q!Lr�rxv[��ǞqB�S��S�g����B��1�F[q�s~��,{|�wuڄ����g�Ǿ&�r�J��af�z��?�k����6�Y�|=Yt���q�~�^k%�M�i�Zݟ8|9��i�7(���'��|~���-B��G;��<���D�N��؅���]�޾�׼#ew�X�O̻HL�8Ҟ�9��xo���_Z������zƯҺ� �P~��_4�8���7��5����������ּ�|i{傓�a�kN[�c{h{'�?g}���J�10r?�k�<a����I��w5�_�Eq�],3�!Gw=+����@���ְ�cx����܇j^�����qޣ��VM�O*}x�5	���1��^}Gm�-nR
 ��[�J1-��f�F�����ꆹ��=���#66.��%�G"�O#+B�������lp+:�͖�$ �\]�8��@e�ыR.~TҺ%�-J
�rk�ה��pI��S-�?q4;�l�MP;k���4�|�湽oX[�J���Z�_�]W̝�a��kZ�����m�=h�z/�}5Wk�߭9+�sA;G<zՁ,!�(J�Q]�-ޞCI��s޹�َ�U-g��}�j[�T��υ�]��� ���	���)`s]��$��ˆ?/s�Z��͊��IQ9'?һ'~V�X|E_�7���IN�s�Em���t�}�%��\�����OV�3��;CU|�?*�?ewԙ��Y�$<��~�:�'��� ��彅�/�vDf�5��:X��$�ApX���w��q���Ia֞}��R8�����]��A!f��ҵ�5'���\�������Iۖ�j��	x/!pAH�Y��Vy Uc��O'5'�k��E����z��+�c�<;b�l�i �� �����o��ɸ$c���xo�4]C�Z�YZI��%�z���?�����q�`���*��glctr�/Ļ��qD��m�,�b�/�!ӵ�*�\*��V��T���k�Ӂ��G?���o�S�^�5Fe^v�pOԏ�Ut7���z~�8���q���.$�F��3^}����5���b���/�^��������ݢy�U�ǂi��1#��:�<׸�Kd�6����ZhD��� �����@f;~VZ��/�����O�����+�/(ԅI䓜W��<a� �����ǎ�MbC��8�/�;qF��$��H�C��>(���W˂%P�@��� �+,��X�v�R�V��������ע�g�𣱱��i�[���rhW�<L�Z �\~�t'��V��n��b0j���A.��,���㚾[l
W>�׵C�=,c�ݫ����6�|-�p�o����^0��y<��q�?�|3�����P�k$o9�v�I�+�������O�����`��e���eX�$������>1h�A���Dm�ҹ?Y�� �c9*�R��6���{��xf�C�!���5�_~#zT�I>��'����Vf�M�*x���� ڑ�~�{ׇV);��u;��ş��޸�KÑ,�8"�A�<��v�Z�b�r{���%��N���G�#V�FUy������G�qZlێ{�p��!��V�s���w��+m5�'
��We�x>��ɤ')#�s-��t�O�]>�q4�[n$�q�]���rԊ�φ�,mW
&����>1|]�Q���w�l�� �|â����Mu^*���ó(���G�j���g+8���=�طB�I�����_�"֭W�s�Ҽ��L�2P�"��-ӧj�_��L��ZH��lZ��ǙU�pf�o�Ooa�⹟�:��3q�F+��%xTG�y^M�h�+�<5qm�4�R\���D\��<�Q�%��C���`��U���	]�7o��ξ�խ�m�� ��ɫE�%Ƕk��i��������Ċ�W��3��#f�x�7��ǭ&�:�3���#��Ú�rx�<��+���]�;��*$��
~�*�\c�k�F��e��pIS�H#\T^-�b�6�,�3c�h�@���v��e@ �s�]�H��޻q�4�t� @8�1ֶ�}�[�j� ɒweg������SIo��)��J��)���A�A�s�^5YZZ��mk���_�Z���i$]͸�5��/�Z%�,�Ƒ�9�^	קM5���k;����&�%~��̫'m�;\�_i�fp��cNo���`����o^E?9�*6�uR���k�����,{N��m:�PR�B�`W�X�?�M[F̓�����:�`�Ff�^���5͋*8bz�u;��U����ܞ����6F��l`��?�u_><j~ �\1��#'����7�ǌnd�n�䌎�WQӠ��x� 	E�����pT�g��<l$yv�!�ۚ�k� �C״�&|*��� � &�g�m
��9H�_.?8es��_���O��Mk&fm�m=	���fy����?6��V�;�Y��2���+�vo.�b�xʚ�m'�/��m���k�j2���}�ڹ=[���u%���I��� U�D#���n��Z���}�6	>����f񕾱�I��8�zS� �S���-��ű���^S��v��%ʲ�'�V3}P���m���Nr*�u i�8$���6�%���>qa^MF���Ϻ}hh�E�UL(�_Z��,2�y��I�a��۵`�;��;)ʱ<~5T�ܬ�̪�NA�C�4�̇ �o�I�i��,ʌ�w��Q�j�?�$.r@#֟k�ʪ8#�ǧz�:Hfc:�l�t�كt�j�I�u��Hi2��pj���\8;���j��n�}(���s֝��� z�}܎?ks���T�Wsdt��Zp^}�7=�t��pT�}��R�,-�ⵧ���=���3���V�%����95��E�Pf�Wp���-l� bO=}Mw�]q�΃�� ���2�9ڼWd�8�$��p�0����hl�\:��Q�lݕ,��+̝/#Ҍ�zt/����
�ϊM{:���4��o������Pco°�o�'�#P�ⶣM��g)���6ڤk8#��c�sS��Ŀr	����?f[�u�e�\� ����5��К��s����9\g?J���8����e�����Tt y���^��*�D��d�m&���t�U����һ��[�;U�2���5�V�.m�S�m��x����7�j���j���,�#a��$Ӧ�"�w�Erzߍ-r�v���S
r��%%c;����J�{��c'�Ez���Mo�T���y��o-��B\�&b2s�f�o�6��K��_1��p�{t�g�X�5�qO�:)@���\��vk�Q��)랝���c��4R���^*+	;3���~�x��7X�<�־��?���뻊���ц�������|u�k������vgv(�>�5��q�y8������}��O�g�yn��K��$��
�='�5݊�'wץ4�G�����3W�V��ȶ�O*������n��C(e���#Z��syd�S�8�^E�x�{��ݵ��4�}ش��i� 
5٭D�x,���n*��� �|ec|�\�ħ9bs�ꗇ>._i6p�H���|n���t���긩��.�<a�^�����H1�<�>.mN��*�d�q�J���>�ℚC�� W��B�5G�ы8_�p��?ʲ���՞�k�d\��mh���j1nnsҸ��
���r�|��A���N�4X�$�N�*������Sr=H�#�-64��.8#�s:�eoTq\��-~��c�L� rf��/��6�$\�܄��Q�GU:�L�c�)�<┯�����p���P�G�l�������M5& � e�����\>�GO�G��0o�����VŔ�mx���i�;,$A�m9����5��s��0N+ҡM�S��ѝ}��?Pw)&��x�5�Ǽ6F+���|A!�e&��U� �Z���J� eM��NG��^�ak\�:��6S_x�'I����q^��=/���,� �}k��1�_i���{)a�N	n?�l�d֦���,��0=�ӆ��Ssk��/��=��e]�+��^D��c�H�O9l~��:?ƭOH��LlQp7�7ǍSyb�� 2�U{>b#S����W���,�s�SC��-��d��k�� �������.9a9��|o�['��p1R��i���K�ߋ�X+F����WG�?�:���\�"���.FO�U�O�����Շn9�i� �h�M�l`��+ rr5�$xb�C�-.x#��<}a�A��iZ埦W�Ep7�:����y�%ws�NkܼM�j>'�L6�u���Gό�v�/m��w�?���RO'�u/[_]�\�:��g�K4�wPI�1��=�x�ٙV�S��יR	���f����\xlmw>����9��[G�4�t�l݈P@�=z�5]ƍ�M�9���� �U�դ��	�3M�
�A� �Swn�,�����969Շ�c��)�֌[���xi^�'e�fP��z��ɧ���ǭxt6^*��-��a],/��mB�H���]�zz3��TT�w�uIq�z晣����e�u�?�����,e�;d l_���ܴm���}8�zФ�c��L��vz��#�r�i��9��<Q�-V�Nj�cy�W�x�?��7��ԑEl��k�u/��iz���ݺ�����^��cϔ�˞(�e��o"�O�ƿÜ]-���k��fҲd�lW��B�6����f��+c�3c?�k������ʻ�ی)��ZX�������+����G�cnx��O��y#���q�]���!�x?P���%�%'��+��1x�kP�x��I��<Qo9P)�Hq�V�i��3d��k6�\�t��Z���$�#�<ӎq���n��[��p�ƨ5�
�ҕ�Ebf��\����|Yr� (��*�
t�2��Y]���Eđ�*ߕ,rK1!U����4h˛��Vw��Uy#�B��ۀ���}YqL�R��UiP��84���4�+�bNc�2�j$��"�#�Qp&8�47�D�I3�w9��M��{��䝼
�d���s���u���\>1Y1LѶ�R�ZزX��J��3��z��Y�.�(���c��;�ҭͽ���;��Ƽ+�?���׼���`V�}6��i�E6� )�uz1�8�I�y��2:�������<T�����j6Ǹ��^��4��S���:?xyWj���g�7s9u<�T��V� ��I�?͇�c��UW�!1)�
zzש\�%�ۛS��U�Z��p5"�؟�Z(�.fv����V6�Y�\ 󬏊_t=j������'����R?'���̮����=*�?m|3fn�mQ�$��h�M%�Жyu���ow4��@���� u����Z��U����W� 	'��w)�.T��sT�<C�[��d]�8f=*���JM�����~���wm���DU9����y���]CÓFw�m���:�y��r>N�_h�\:\��e?	~Ϛ���f�g^�̠~����E�lD�Nߔ�l���7�-Q��˞q��湟�����e�cw8<�����r�Z�@��q���� ֦��#�ǵ8n+�����IL�C�AK�{�H��Y��E!�~�V2��ݏ�)m���~��w���a��w0�k�//�I���?�|!�� m\����yY~���{P��y̝��=�@�i9j�RF��ԓ���m�Ȥ��4��^Mԑfh�����������E�0n�����n�R��]ϸ`W�~�T��b�tP�8�x����5�\�C}'��]h��hI���ܧ�W=MΚgEqo|;;xO[���O�jd�o��N�� ��_i�q<�y���� ����7AG��1R=	�r�[�Υ��]􋅷�s�֫\x~�u��C��e�&x�I	p���GJW���Hē<�yg�~����G�;���\��c<�f_���袷�� �q?�W���=nf
oZ1�0�I}�{Y��Ԓ�O���P�D^ѣ����\;;"G�#�Z��,�"�(�{�����ŏ74�3��v~��׍�<�[xeLϷ�J=�\�g��u��a\�Fx5f}?[�@��P>�`�ּ�Y�������;���n�=Eaj���7G����u(;��O܋�3�Eh���>T�N����_8�y����B�"��Ǧ3W>�`Ԯ5D�iL��'y9��:j�P�'�L���z=i��4ϻjeݾ�&�O�!�'�b�B�&V��V���6�Ma&�5���Fq��]�����$�������쌔Q��~��%��^�AԌ���T��5�&��$�k�Ns�֟�/mis���I��� �?ֻ_|`�V���A���s�g.e�Zt>n������ ��p�V۹<W��khd�2� �۟�c&��K�6䟽�Ӛ�e`�M�U���yғ�Ҿ��]�-�/g3<I��`�z��_ �OT6��#/#7�J�c����a�����}���t��+)n]�S��Ե�!�&��?�e�ƺˇ���OQ����x��Z���e%��[h
�� =��׼?�7�vv����}kg2e�
��V2�iٳnV�u�}oc��#�Qӹ�bry�n�*�9�8�|��5��f��i|g5qu/Js4���k1�CK��+�G�I���HE��f^�����6���}��9����&��~�>鿊�u�mVhv�ܛ�_����<�=�-�rn�Q��U�t���*;����F~��U����)�Hs��5���Gǚ���B��@�MG-8�ʳ�=���ƙs�F�����[K���	u��q����Mx���6��W������x�k\~��-�&�$�B��JC��������r�}�ٵ��G��4��jQ�9��5࿴U��z�0�.A_c\�j�?������.�5�|t[�]�[*0w^��rkhǪ3�ٙ�?���YWp�{��[�T�gr�mn���ٮ� �1)�x��d���j�~�r��#W\㺑�z�5\�B���όڦ�g囷`;n�u�.�5Iu+�$�Kz׽X���\*�����?�yo�?�� ���/1(z�����G��(N8�o3�?Z�pʢ�x8Q\u��T��\�~�iq�Fn�d� ���?�tY4q�XG��h���tw�u	��z����{5�w��z�+S��)��,xf���}�3�H_q]7���SD�$�F������>�.������+[ᾭyd�#-��iJ/����{/�����0���d69��?�a>",&L���J��{���i�0�`׊�y1�N�+u���s�_
�wD�ɋl��'"����t�TI"I�H<T~�N�������@կogl��_j�q���%m���^�qx�5�V����{��c�&���,6(Q��f��v�����A�+Ц�5{�y�S��(�/=�Z;�4�#��� m=1\�2H�6�Ol
�C%���~e�����}6�9e@�pFkݧEYT����|���R%�@F��U���ֺ�ĮK�ۂx�SᗊWVd�#*������sN׾)�>������� Yr3��[IJ
������㿊ZH��#�����ʽzZ�.�b�[I��]��~G�_~�������]�Q�o?,J� �,G�^w�|P�����Le��y2�Z���O�<3� ����L�ѻ+���Ǌ�߆���"�܎�� �_��+��6�0��ҾJ���i��gTK6᎜��+z�)��Bg�|��C^��t�ž�d�vz����.�<"�K33#e�5��=�"��S�H�H��t�n���ז�7��Nzת���:]�����c�W�V��d��o�W����W�K�����Ky�O�������]G�S����Sm�x痐�g W�^9��c���z��PEyu��[�iF��.��)��#:�	��M��]W�?��zΗ��5�mrK�U�cT8��ֽ���"��<ٶ�~�"������5O�:����q��#��y鎝q�YF�IJɔ��(�t�,u	x�;	KI6��W��P/�`bw9L���Cč��R��8��昝���?ϵu� <��tR9��${׵N�O2��dx)?�;G9�HO�e)#(�F���WY�Üb�C�R:T+R���h$M�[>\�L���p{c��Y�ju��O�/H�h�`�?ʾ�����9�#_v��&:,�/U<�¿!	���ɼ�����b��	���W�"\M�D#��W�<-c���ݎ��'��5��p�3��>+]\h��D�,bO~��+���V6uO�z%݋�����>\q^?��V�NՅ����7g�z_�f֮
��ȸ�wqSx�M�,7h�3��R��>T^�� iiw��ҳ.�e 
�����D�h��u���W�U�;�ƺF�B9�q��q��Y[P�h#�������U���[�~%�H�o�s�z�O�sF�C�����<��\Z	X�3 ��U_��,6�	lƟ(�{Tɩ+�fd��v>��~� ��ۜ$P1!Kg�����|	q�A[�!b�`J���k�I���	0v�(rG�j�/x��\�f�V�,�x��V��j;��c�Ą�0x=sT5_�^HLw���oMh�A��rÝÓ\v���q,��ݔ'嗑����ȔP鵟�Oٕ��6����O��o�d�;���g5�ç�{V�w��bvV�,c ��_
x~	`x���/�a�c���]٘�4pV�2�0Qg�����Wg�jKy��ևdX$8��}���s.�ָ+,^?A�Y�d���(��1YJm��(���\���0o�/��|�d6J�����τ$�]������-���>�������u;k${�q��@�����E��fV0�Ьx�N1M��'m��3w���y`�#���'$c=+w����Z"�Xm��|L�,*w�^zV����2�v�?�{q�y�w+|����e�C/?5v?��}^wm?�@�^1�^�j��݉� 7M��5/�z���7�T$V�����jM��Ipzb�w�͍���u"�:�~ޕ��c�F�sX�ORqV!�,��0!�`:)K�V�Gs��ӭ��Z����/�*��*%?/�Z/o��oGbǠ�q�]�����6ߩ�xf���V����m�c����֝s��`�}ˠ
  sۑ_=�.�	u�t�P�Xu�����	<lbE��x��D�)n�I�,�xS^�տ��P�`C��9�__�n�����f���N�}��\ x��wÿ]i"%Y
�7 ��#�x��sɝ��¼*��=T����x:�[���q�q)$*�������?�����z�����ʔ��י|mQ6���Ƕk8T��5�SG�����%�S�ק�jh��%��ź��Q� 
�O
�i~�3Ed��v��ߊ��>=��D�P��;��^F�'�h���B5��T�s^��/�x��D�tcoA��W�� ��L�Ʊ�0�(�z��]Am�[����c99j�#����~񕴗��r�w�}_�������@�#o��8����E�3��K�c7/=��5�n��ۆ�y4BҒ������6����5E�.G����W���,dD1�GS\��V3�WE��Ew�<�,�����T��3�+ކ�<�nO�#ĺ��t$���ug㧌56��ȸ�	��K���<7��.k5��P21�p�Q�oP�m'�ر����J�$�~�J�d�H7�p�����٪}�V}� b���4χ��k���{�9$8��+�>7j6�z��"����kVGS�#�S��O|*�z�/LQ����eu�{��j��I�s�{���rX���B��=+�4�n7/���^��I{yl�	T��بަ��E��<���&�20��z}+��kk����W/��6X��I������w�{K-)6]�(���q�w���K�  �tZ�K{5�ԕB��+�<E��u�NC�~^k��x|�P���ݪiE82�7̑����M"-�W�^o�.�;[��s����{�p�[+}=+��������`�<}�£�G|1�����sֽcP��&uix�Z��Eoo�F��<���Ko3o<���~��|�l7,�@�n�����İݸ�NzԃT}�����d�<)��tz��k�ٕ"��9����,�'�7�[sN�G��x�0~���V�� oH��!��zS�I�|�=�����8dA+l�6�V�5fO�^]�J8�#�y����ʒ�bN��������p���#�"�*�R���.ō/���{3��������x��T��0Fk�-�ج.R��H������f��ʃڷ��R��H�7���6�ӿ�u?u�<;v��q�Z�� �ߗ�w�I&�>#_,��B=�z�Z���ǀ>%O�ݘ���g��I�>+_]B��>��'��=s�f�_R|?�t�N�Lʳds�W�Zj2;�a��L���sg�� *�LW��]�"�y�#��h���M��*�$`VW�4�O��Xb�x��cN�,�%mO���uo�Ii$���S�]����+� 7�y���G����mV��^�����NT�<��^�9sX�+13��������C�)\{��<�"�jHۏƢ�׊�?�=)��p�7���4Q7PA���:��'跌B���i�>"u�����u���c/�K�8?ʾ���u�p07ʼ|���b���L>f�IF q�^��/���&Q�Ⱦk	8ȯ�;�E�_�������W���~�q�a��g����zƝ����4���Nw
��ž$�R��y�y�|W��K�>�%���X�c��'�����w67l3�i�N;�).����oxr��Bj�(#� �]w��:j���6���o�~_皃�2h�$��������]���� ���)~�Y���L���B|Oզ�[S7˸�v�_H�x%��p9�W;�;�+�k����b6 �� �]���w�.B�X�y��l�`����w���l��:b�1��#�8�0Ey���[\2D�hp����A�?8�5�Λm��d�{~��v��=A����P���� (j��Y��� ���۞{�\���9t;���+n�	#��aӱM�=�v7���5����g�R	� 9�J����;�"�1�; ����z��k���Щ��~\ 1Ke�����7IQŎ�� ��G�������ܛ�k���l��?
�����1�+�5Z���L�ݟ!}=���.�Cd�_��h�Gz�Qi�h�:+�j+�=2xϵ-狡Դ�������%񥼗M�8c��+o4�2/�H=�[S��3��:�����-9��{�U�aeR3\��Co�-I� Y��$�ֽ/�#�E��ې[�Nk؏Dy�78?��*�a�f&�+�^�q���a�lWܣ?�z�_���O�"�B�?J�?����+�U��I��>Z�>�R���3�L��Ś�[,b@@�}+矌?	[K�[�5C*�с�ץY� jx/�)ڴa9��j���M'����V�y�,�@�s��%kyp�8<�Z˫�7J��%xG�7R�HT"�}+��4�qֶCiI��ЮMƯV��+�X�� ,���a�~� Z��ñ���0�d�������u�t7/�b�����Q�5����$W~^N�8�+��ܞ\d��k���#��]�n	=Y��7���O5�T�wsԋG��=�7qI*�
�+�>.��⨉,T�K�����m���1�s�q\�osVf�yeO�;�"���m̏��|6� ����	Xc~���^(�/�5�}��.����`��+������[ڭ�kgn�[����G"�y+�d�r�g���E9V3!�<�ש��֋$��}?�U���6��5���s�#�o�S�}+I�Z	�#
sS+��_�I!�$f;T-�+u�hٷ�u��8�7דK��Ǣ��� �����k��-��9t;o\Gq�067I��5�|g�F������G�
�?��eǋ-V���������о/��k�ޑ�m���8��ڎ����x���_x�8�	��ұU�d�Q7�� �>�&Gڧ!b�6?ȯWվ#[xa�����@���T������\�(��Y6>.����ڻZ_�+I�]؜�+ɵ;��B\�5��ƿ���5֝��K�|�qi>�t�\�h�̧�i]�f�3��P�`f���OZ`hh��;F=Mw�_��>P��^���[�jH�N��d��y�0�O��nUcoŚ�j��e<��� ��-=UߐI��^,����m>�������<?2HJ���cѮ��}:h��� �==�_y�{֋]H��'v9�i
�z��a�W)_Y���z^��GfT�����ڠ�h�yaިEy�
�@��]�eG8ȫ��܉bUM��Gk� �uM�%՜��<W5�� �Z���6�b��&c��{ק�����z�D�+�����9s��.S��)\HÁ�ޢX���nM{� �3ރ2I��lq���s����i�<w��Q³�ֻ#��9'��������X�5�c�+�K�6t�v?ma��8ظV#w���f�YՏ#�&��˥��O��ܶ�,j�m<�x�d-�cP���l2��� ���Lt���V���4�������d`=�yG��]��p���<t�6���-�'�� J�[�Vj\����m۲G˓]���xGʊ[� �\��y��G�:q]o��&�v������ ������\<:�w��_GxŧL�Q�"�m�Զ�7`|ٯt��)�s���1U9Y�т��?��fa���<Yի���1\��ZNW�Tsm[v
>Z�#U��*:]��&� |}��5��괞���^_�>����~�� �V��/��A���*��<���m�*�da�ޝ���Ǡ�����/�^����p:R��#֘	�ƿ6�sA#�!2ǧSnF����:��'���~pJ
�C�&[Z����}���C�~bB�~5�o�L�zr��b����c��lchW&�b��ޛ}y%��d�c�U�`�ׯ_j3�^��ܽg{$d��q�5V{�g��9۟Z����}�8�{�+�v����F��+Z�x��G� x��`5�\g4n�b����k��37w��,���O�حn.�#�Ilv��t{?�jP�lq_Rh����:)�L���&��4�>� �}���ԥ�}�l�VQ��P_~�z<E��9�-���m3�^	�ID�3H����P��K�4��[���@?�\�-�
o��� ��$��\<E7���ѫcTm�c�v�D�M��<����O7�L��p*j�#Q�u��\p5�<�����O�:芻�X�(o� ]w�7��u3H�;�� ��3[��"�~QX�6>��
^ėP���g��Ӫ�o��V���[��ڊ��p���_��l��bӚX�χq��������*���o	2�ט pw�V�O�b��w��.73]�)�o �3��٪Rx����!��2+�9�i�m^�S�T���s,g#q��:�/�������
���	�W���"�!�rH��^o�EXir]$��rGմ/�sN��_Vm'RI�o�@�^��t0�h���$����m��=kFD\q��qRј�8�=7�WŇ������:W)��ˣ�	�ڹI�3HI�ڒ3��8��V�!˩�x��\���`WW���O�Bϸ�Y����zT膯=��6l����φ�|9�x>+K�0�TRyǵ|ţ��Q��C_[�&����<2Mh���� <�O5�Chhq����ǜ	9���j6�s�S P�s�-޵������a=��"�����H��U#�ι�|��fc�>�E?�j��ÿJ�J�)���um��G��7x��X�g�U)~.x"E9Ҧ+� \������AT��G���l2��q��L�<l���� ��[���&����:�0���|l��B���0?�/e�͜���|;5��A�1��+�ȸ�&�A�T��t�cH\���T���������+��v��Rw4�{6o����VB�?�ǃ��������jWnJ�|�ƹۯ��,q�;��+��5J����!U_��'=U����5q9_c�|-��i�#��<� ��\��O������PS��|s�5K���*F�� 	�~�ڥ�\��F�|g c�[�.�=J� <���{_�w��,O�?�~�<�Qõ��Ő�F"����ĉ俅d�ʃn=���������%�O�2���m�N�	ͭ�����JW0#<ׅ�\�s���O4vR:7B�s^��� څ���[B��͌S�O�B�{�l�D��q���(�Ѽ/����� �qJ�ץ?&�s/�����m����`�H��U��\~�1��*��#���~��.T���ԑx/�I�˸�� `��������fF>���@@�� �r�1�ƕ��w�<����\���p*տ����g�]��O,��W����)�Q�l`Է��m����(��Fs��I<%����2�?t��+�#�5��� Z��C�����@/�wF�x�;��!����[3��_���r����������߼��M��b���X�<��h�6Ҧ�����|a�K"�ǿB��s��"���rх��2oFD���=O����� ��P%?>~����o|@���d�KnW#�5��-�E��nl�[b�)��vW�<9�`�r��C�RN?�)�r��s�h|a{&S�|��8���n.�o2|�:g�z����f����Lz	O_��:��xt>YΧ��dG>�)&W��~�'��NX�W=�v���gs�� ���>ڋ-_�vR�q�z����Mc�,�>u�3ҹ��loCtY�k�CO),���+��^��t�8��sy���>�ף���8ZFa�Qɯ��;�g�з(����|D�&�,�`U��N��>�2����k�p�Ab���}1�}�L�T,O���|3�t������?�+��E�.�t2z�}Z��wse��4�r�9��]W���;�6cn���Ҿ�G�u<;E�����0�0��������>��;��nf��؍��z.��������v篅z��#����v�*�xS� �@�5V����W�ӎw.+ˍ���JZC�h�kH�������.��O(�T�y���ֶ�~MÎ��3+x<4`�(��_i��Q�ح�����������?5)"�U���p��ղ��0�J|^�d�$qo�o>�R
��T�?D|X��(����?�B�֦������~(C��r�3�W���'���z}k��lz�����k�X�B�x���M�9�R�+l#xQ���\k��p�k�/x����p��k���Nn.��k���S��t�v�{\�����9��9��������/f�kub˃�Ҽ�����������������(�<ݙFOA�S�i���2��I0$��O���u븢�Y��7aO5������wb"o�2�yw�:�"�3��!$��#��G�_J����X�w�[��0�~5�ʀ��`�k�g��S�����Jʣ��6�u<�����|s�si��ɧچ̳7-�N ��+���M]'ᖑ��6W����]	$(��|��w�W^�մv�\"���
X>�����h-N��P����Qc
�H'Z���jZ3��q���֞����{���,�q�ה��ᆐ�3��,�2v�7J�6�R����$��s_?x���zF�:�p�ۏ
z������5��W!674\xO\�2')��#��v���[��ź�"KK[�Ш!�6o�Rjx�<��}���1�]X�Z�{�u��ۻ����5�h� �HYe�I%�O̪��^g�W��"�Y"�r\��^�����X��ۙ�� �ʥfތ�4����ᇀ<d�]����.'���5���g���CY���C��v���Ǡny��x_��%��@h�eU=ȯ�W��`�C$b�D�W
�8���Y�ʹ���b���� K��H��hیz�W�G��%�0n��g��Ʀ�gs7V$���_�{t�bIf�S�sͭ���%�`u۟Zd��|���F{ъ�I-�X� �4dzUhHҧ[Kf��A5^�1Pj}JM��zk,����g�q���'>���_5�|jP��k���k��r�!R��G�X�:)�q����� ��d�l��j�b��`���$��1�_T|K��|#�����Ŕj3l�G s�_9|	���^ �h[�u�[x<�5�~,j3Z��t�$-��w��䧣=��4���jm=�����X@
x�n����+Ú���]1�8X\����D�H�؜���^K�[w�)��M��[>f��O�S�����HI�4r.�t�A��(
7A�S.>��Kv�M��ߩ�� ^����뷌>�cM����Ǩ���*Kr{��>���A�@FH��M�tm=��♔c-��z��{��z6s��g�v��m�J�w���Ք�>��I�3�~
�:F����Es�J�c3��g����?��S�������]t]�[��m���#־1�+��-�w6zsڽ�X��u�$���2�n�� �Bnm6ʔU=���[/������@jV�(e�: ?Þ�����n�m���q�jS�����C/��k������� �2�Rkۅ�H�jIs]�Ue�_�>X'p��Z� -����g!r��p@>n����SK���+0;�W�˘l|a������X��;�*7`��Gӟ���K��h�z�����̆�&W}��
�h�w���}Eh�"6m�1�ں� �?-�t	'�X�98㎞���!O�^kh_%�q�MxNsR��S�l|�&�o&������p3V|D���5E	���W�i俵\��s\ϊ~��(ĥ�Y�Z%�����g�=��Ĩ!i��1�wҽ2
E����E�}���ǥc��#�`�8X�4A�`���֍����<�d�Rxֻ�	�N��%?�c���־��~�*�ï��(��
XK�0�qƹ���E��g��'X�jv�/˵��>������mV}&�+V�B�5���>�&��˥��F�b�+�����ԴKI��N{�1[ѓ��f⢃��C�Όy>����W%O>a�u�߳��H��͸c
���5��b��?]*��HH�q^�>r��<?�k�m�@�
y`�?Z۳�n����t�"�C�:%ƹ���c�^�zz��C�ߊ���v"A���A�3W��ɖ�k�k�{Y�!s�Mc����Im~ҩ^0�+Ծ�ĺ^��͙���e�����kk�
���Vu\�i9F�Agc翇�*�A����5��z�h!#�����N��?$l��ҫ�^�Hu$m��Q�笎�;��]qok$M2���&���K8 �UI� �+�m.��B2� @�WQ�%�UY�q��x3��+��cQ�I���\+*9���o�^$�T�,�A�����L���#��K�l�XȲ?I�]��&�k��;��z�������WT�Ι�ʓ>��'�-����n��� �]�����!<W�s���h�h6F�py����Ml�^E|�-�/Mv��'��R|�+̭O�G�JJ+s�ˉP� �a�W��Elr1�Z���"�Eݼ/Кy�����M���0��6u48/*I�3���/"��a�myg�.��ZR����z���_�y���z���G����y�3�Q���}�~��H=���+�G�-ħǟZkS��Nis.�G;F��'�v�EI���oI�K�〹9���*n�ܟ?�5�7����8,G�k�ϊ�n�'=N�+���g��'�Cx���Y]͞>�������"��DU��\��k�����1�����[���l������Z#�*��=���:���v�m����8��1=���ز��9��q�|Qi�M%�llW/Ҿ\����v> �n� +x�J7����)��
d𕾔�;A���G&���)�\Z�}�E
z�=��=a��إ��8�z��I%�Ļ�����(���;L��"�o�e}�/�����Y~9T,>ּ�����b�b��^�i�:�+b�χ�ns��%���Y���R�� W�C�-�R:�!�#9���êJYv�rX�߱�eP6A5�֌��=�ZǪX�\�O�O����Ͼ%	?�YdUu�s�^��=Q��۹���W�x�o�%��w���X�4h�������F|#o*A��Ҧ�ć�b���9
w.=y����<C�;k�^;�0�A�Z�toG{,Z�]B~b �B���3�>|��_�I$Q�o3�F2y�{g�>��d�?
�'�$L���rF{׮�6Ԃ�0<�'ډ_���W;KZ���vt�)גM��	ER �ך�/x��n��s��n��s̮Zf*
��c��Q�Sү3�|��[?λ���ɤ�V�kɴ}i?�$�L1-&�޽'�v�<�]�K(�1�{���+@�76x��i��1�3Eu6�F6�uR�*)V�d�sy7hq�7@?ϭ}+ky%�����P�z������)|�d�'I������_/a�O�M��G�xkZ6:�����k������9>��W��Rb��Mtv�*�n8�t�x����S�Sؼ��c� F{��1����H'�=�1Rx��'�2�9♡�o�x�� ̽Kt%���sB.��l�g]��I�q/��8���c>����>D^Snbs���4�ú��j�,���P�N;V����.������d?
���2<�g��`��n�e�3��p�5�����$��5C��|7x�G����!20V�g�C���lfWU8�Y�]�ce��������nq�����P\Cq,�q����y��Tl��&�᳏¸��yu)���ִ�գ*�����������Ͽ��]��I��ݳH:���y��M�X�`N�^��SO�Fm ua��b�x�d���3Լ�������U}����uҮ�8�R����G�6�s&��!w�[� ,^��;0۞i��2��)ji�,`�nFWh$���y�G/�~�$�1\��[CjG;� �-������	��xRL�����&��L��[���y��c �>���z�����Q�Z��E~&��8�םZZjwS)��N��=i� �2����+5�ɥ�u�9�:-P��qm�6�z���g��h�ye<{b�J��נ�]}���j��~�95��K���1t�B+z�I$��8�5�-`j*�p��xϯ�+�Z�������pՕ�OI��b��k٢�<�3ҿg�5�r}?#\��Ğ-��w��n���������F;W7�~���O9f26�I�Z�<���
uY4�O4;U�3sָ�[�6�o~�0��aX����|Yu���M� @�q}%����=8�V����ǧ���sn�rv�?�Z��=[^Қ��
F1��A3*�9 �N�c`/j9������K�(���2z�W�6Z��axTx�X~���DKl��>�����o[���+�3�
�Q�Έ�����d����9��6�#6A��k�i</�	���w�6�%��j?�5M���J��U��J��o���0������|��]�9^j�]|#��3�=& z� �v��kuVS�q撇[�jp�|4����(*����+�<I�k=� 2+6	�j;�CE��h�W!	���v���T��M�:vWnޕ��+ld�|�X�Y�<�dv�>���3۶�6I�c�+��C�2q�)n�FiF��)!޺L�� L��:z�h��2� n\@�L�ch<Կ�w��Y�ORk�h|;�X3xrX�Un������h���Z=�a�c�X�.�(�&����H9��&�ܖ~zm� J���[H�g��$Y�����1�:���E�����>\l6�kXŦaRI��&O�?֌c�5��f`�� :S�Wb8�E=I\��v���M��f�$_�qE#��"o2�q�21_|T��'���}��5��=�ʾ,��n����S�ۜW����������=i�}U s����ƿ.5�9;y��O)��4�$2JX��l�͝߆|y�BDRQ����O��Yp�1�r��c>��3n&�kqs67��Wy����x~��)��k��~���C6��h��{lm�x���Z\ ݿ9?Z�/s\�-ź�ѷ���m��gW��$W�x7�����m$K,c���?J�q���.�������>�ц8�9?J�iu����$W���<!�B^��U��
A��c���,� � v�YSo�֪��]7�Z����R���3\�����4���?*�+�|c�������������}�U��ؾ��>bi��&�nF���5z��^���=̋��5��焑r-��䆚�<#���\�
�G��c7U^���@֮$2}���8ݴ�]����L�H��(
1k�����7l%�|��M�Oƣ��o�3Q�iob��<Vm{T�a���� ʗþ Uf6s���b��_����2��#ҕ�2xus�<���5ҩ;la)��� ����ݼ��yj�%���^��z�[}�z�]�w�k���բ�<�5ݞ�c���6���6��R,P!
��海I)5�=��ǵ9��$p)����(�i+�)�V�Z=�_A�n��
�C�{6+���G��a���9�4Ql��hD�p��?�}A��K��=�;d�!C����� ��=s±������H��ס�?�Ⱥ�����0y����-�����ÿ6�>4وsú�mAÿ�
XM��k�����4�S�v9���0E��4si�6��mq�]�~��C����>T��ƽ6�#y�Z�gM�oː+�mG�V�0�U�Np�g7��y]0d��@T�6�Ín��3��t�w�:�K׶��-�U�`���}���w����� ���:�,�m}1Si��G�G�mhӹ����L������MK��J�Z��T��W�M�oO�������ni� �ȷ��� ֧�X�ek#�n�_ȮZ���tlq�w�m|3���z}�oP���^��-����G�@�M� ��l����Z=�D���k�O���ZG{9�RA,�@�kԾ+iw����<gߊ���H�#U �?.Es>%��K� ���70��o�X@N���ǽu�7�j�,�����' יh�����/������;Ao��(�`*�-�����ټ��� ��;����)����n�v����5�M��^m���R��xa�H��F+�XyQ�;F�&�k����B@ǥQ�<A{$�ƛr��i#�V��e�.ŴEq�Z���~X"�5l`d��ןS)Q���`~�?��\)��6�{�l��g,0k��e�<Y�����A�]H�\�Z�9#i=�k��5��b�x�ֵ5��6n�
ڏ\��-Lqi�{�8�/x�T���%�I�ƶ<#�k�,Q4q�inO%���L0n�S9b�<o\𿉵+�o��:�r�ϵ2�᧊.Q1�����o�}?�v�����q�ӊ��g�k~�]f<2�����SiX�CG���O�6�K���r��^g��HD��Ēz
Տ�&�*��W��J��jr�ڛ�#���m:n;�U&���_����lv���Ayϥ&�KҌ��x"�4�����6K;Oj�l��nx&s�	�:�%�4���Z|�W��x���fa�0ɪM�O�M��`H�>8��ᔺ�򫞽����[9�W���Rh�R�G�Z�=b�[��h��
+�������ul-�o���wz���Vb�	&�;��(�4Hq� ���J��r��H�&I�oLg�QI��ёX��SV���L��砭�{����C�R�k���c������V��e��mml�m�@�s_T^A$ � ��N��t�ZM�#y!���KS�dz?����#��oZ�Q|I��j�T`���_4=�VW��/5�_�?G���]ű$�~3�T�r�}��t-BHU���JĖ�^X8���|.�銾F�\R��s[D�oP�'=h=iOSI�Us!=i���oZ8�E�+�g&�l�'qEI�6?B�%Ŕ���ھ1���^��I�}���Z�A�1���u�1��� �^	�Ǳ�^��q��:���S�5�
3�<�f� V�)q�&��`b�^]J�B�>�-�9�"��^[�"��u�hŗ�Ռ���Vv4>����$�9�;�3�����Y�1�y����B4>�� p�id�;�y�sֱgYx*=jX]��i�W���oُ�4��K�K�w�w�7�zw'���ѝ٧Gs�?J���I�(�7e�o�:O�s���ޜQ��M8u��T��k���T4PEP�N�j/PM3����@�n}����A��a*g=��^�V�m�)#W?���A�������|�:�?*���x��R\�؎�a����W�z���?��Rf�YT�F�z���>�⦷��-��;W�q�5���5q��K\���1Ҽ?[�T�kS<�U�ҍ��m�})�?H����ki#s��s׊���Ǘ���?�Б]W���5�~�7�6�V�ϊ@M����#i
R�lq�^K.���^����j3G�j��G��8ǽp[Q�B�g��M}U���]t���t(���UVn�AN:^�MR�L_��l��%��~U��1�Q|�9��_d��{�&���Tc"59&�b���Mƭ)��@T��5�6ʚ8���s� �U�Մ<+d��R���_-3�k�����O�E.&����Z���1Ң�s�R��`KZ�Z�#d��{�*v�"	���!�:ʾ��Z��>�+ʖ-��Vǚ� gܪ�N*����l�f u���խ�e�:�T�� ay�*c�w-���-Ė�F\z��:��(���9��zp��n���i��}�)�F� �@�i���Ǔ8'�Y֗��=M^��5�FWW<�?�  ��l�Z��J1q���n��$b���=��Y�v;��;ON� ?�)^ƑN���i4]���� {
�7�*��w2LXv,k�����-�z`}+�.v]3���cҲ�M]�I����bX��c?(�4߉Z�btX�{� מ�]y�9�;L��ԧ[Kt,Ҷ�qҵ�!JW;}3����0I �C�1��\�f���觻��̠�� �R�?��;��2�W��{w���\��_�/��Mr�r� �^��4�]�ax���EC�{U6m�I�Q�gb��Ӊ���op���o�H��׊\u��[ڦ�Ԏ�x����G�ڮxz�GW���e�GjM�i�����V׼ ����2�9lq^>�^��}Y���m��6�Z����8ⶉQ#�j�Lv�+��o��K�]�lqY_M������o&��w?I�?#ע�E��H^y�W׼i=�ݼ�G�@ t�G���ڎ��P�לw�Q�)$���t��14��l��N��lsu;߄�z�������77J������������ ��\���`|?}Nk�n<_m���̨Kq�±w���I8�בY̲̻�s���=��Դ��#�������m^�W=��3i�}�a�<W��7��Fe��<^㜊�%e`���4����9�9�ֿ�� jH@{V@�_´G<��iiZU��V�9Wh���y��(�go�)�ܾ�R5����6I�+�o�V2.�,�/ɟ��
��f������R��t��I(�S��F�g�p�q�֞�O��n��ԩS�j�;����W���^,��O<�)���!�٧���B�>�)BdR`7p�@�22?*M�1��$�\0H��T7ʊK��Y�z���H�a��ԑxz�h�2�����C��/����������b3�������Ҫ�!���Iq�c�W��Ǖ�ڑ�\���Ç��-��޹�=��xf�Wp`O�f꫚�-�5B��Q�9�qPI��<��}�#h�k�����@�zg�?0P��,+��j��"��法x�cX�rD^dm�j}:Uk�2�͹\�[{��j�5��7|{QOU�8�Z��Ͼ)`bf\A�I��2Ӱ�>��_�I�xF�]˻=8�����Z�'�l݂=��4����ӧ��#GzŎ�Sr$f�5����D}S���o�C2�ۜ�z��o��JMY��M�� 0<]�0�����*��N��{�;�;99��c�O2�=O�?ýv��ιM��?�d�N�s�ͫM:@
��W�����@E1�cPk?��������M;�Ovǐ�Y�i�\�Q��垬�$��� �gkĚ��<�9�x���9#ѧS+�Ϡ��I��$�������I�6y鞼֞��[�]>�5�����#�MkVD��nݫ�~�f�|���3�ź�\]D^�6�z�D�]��cI�(��x>-+F�l|��ֽ}�U�c򯛭'9j{t�ȎP��8E#�\v��Őٟ�{�峟�YZ�����s��u's�w��s��6�|��K.?
�~�ñȬ]s޹�S±�q��9l5�x���аܜ�Rj����ǔ=�^�&�-�p3V�L'#q���fe4�����4K�\�����	�P��k�2�!0:�ה[���W�a�9$x��b����lx^�4�F'}���J�p�l��+r��n�8��>��U|m��kt�+���k����r��q��,��s������eucj#Y
�qҬ���F�H{�<�7+V��2F���'H�t��#VQ�m�t��eo�vY�����^;�jR]���%��5��_j6
Ds�Q�q��|����r�߄u�i�Ю�4n
��ڼ��?�-.&��;�3����q�+U���g��ּ]}�[�[�|��#!JWG"ѵ�n�Ԕ���㟭;h��9�yd��3,Y,�R�N#��� s� ֨-���G% ;�eR���:nb5�d����7j�_�/%�7֩M�!�A�\��u<5����}�´�=s��,�����{s۶���H$���U�k��+jsƜ��>�������KYÂ�W3���4�T]�{v��꺥���ӷ��@��� �^ݓ�R��_n����%k���5(X���"1��}j��?*�°�0Tp>��ڦ�{my\��56�⋽CI[}��t�:V��h�yE�s�ΰ� ��:��;U�?ó^�I��5j���o����Y�R�W��p��|7��H�]O�<H�7q�傞A5�]irZ*����T1ܴ,�+X�S]�eM�g��~�m�?���s�J���g�i�Oo)O1wrzW��7�.4�X�u���*��F����n5q�z�}S�ш��W9 f�ՍJ�n.���3�U����c�n�Gw�1Kʎ�R4ȸ$�������НDl���.��P�Q0�N1�QIx��G4��vo�ap�p2qҊ�>�5�~ jr0�H�����t���b#X�F\�p7��v�\�� �kYC�aӚ(��������⥤6z�c�y�\�r1=h����ǁY+�i���V�034y��ڊ(�c��Z���Vgu���MWm��:W;xSi;y�������1��c�������)��C��x?SE�/��GKn���1L�c�آ���w=8��ak�#)%F}k���e��z�Ezo���|G[��ċ�j8�e�v��Q^MF�z4ֆ}�(�w(5��(���QEzXs���lr��qO264Q^�O=�5e~��<ϸ��QT>����	���ޢ��D�[�Ge �<z�Uh&x�r�UK��L[�3��qEL]�1�r{�ϼ�4QR�"�<Z�=�Y���G���l��� >��J��7#'nk���(��������Ze�ފ(-��^;��#\�QR3�ԑK7V%[�R[	�=��b�v��� [���4Q^�c�������c�ފ+�<�Uk�;\�O9��y����#i���5-���k��QP��\HX��4�2f�+R���JҸ��4Q@�,?y8�
�-&�8�Ъ%J(�ݎ�?�Zt^x��
H�2�6�+͋g�-�GZ�fZ���H��	���*]/ⳢبQ�QN���21E瞙��[ƨp��谣O������|�/�#��$X�
@Ⱦq�W�-�elg�F��+��E�Q^�c���e>�*u�����Ez���d31��h���S�Tv#���Px�4���4QJm��-HE̥���<�^���B��<Gmպ�FU���ᜟsk#�?��%����Gmi�c
��EW�-�J;��PK   T�T_��jOw  � /   images/cbe86463-f5ee-4cb1-a8cd-cff047d8f75f.jpg�w\S��.Ů(*(
ֈ���"&�W����4�cAl("RTv�Q�)6PEDŊ
�pѷ|�߹��{�=�s�9,���k�Yk���O���}��0��'�NNN�%}?���Φ� 4`6  Ї���u ���Ө+}���ê~U��q���p����v�O��i"`�o��4�<�i�_>}�� sqw����}8x��������Ֆ�~������7���k ���^����������������4�R+�Y�>�
�I烓(M�8x.x.�@�B0$@���R  Ri����jH�V��s�@�Ph0E���A��(  �*�o�3V�j�?8v������  ������0H���Jh�)���>u�ߪklv��?87u�?8/���~�8ҝ C��=�>��.�;�S_�����>����A���t��Ĝ>�/<����ez��\��P@zڿp��s��=N�Qx{�Ge�q����3�o�7��	��a��9:��P���'��~~]�\�a���t���~R_�����/<�_x���`����\�o�ۇG�G��jӯJ����������w7�?`f~��{I��r��p�W�C`0��T ���{��U����e��U� 8� ܼ~��T�?J����hb��X�#i�q"�\R�� s�`�>��[����[c��#��?�� ܯz�����/��Wtk��}����
��@������8 `���a}�o55��CQ��W��?�A��O��kl~��W9���W����3J��u��9N�O4�����Nk�q�����.���w����	 0x� �A���2x�p�Ç�9f�(����L�����?w���?/��A��!p8�{*	��Cu�4dȐ�Æ{����5���z� �
�Դ�T� 7'g7���w_��~�?3d����A�����P�w�����8�җ���_o<\���
A���ܡ	i{�aN^Ǻ���j���<<'N�>c���@D���	D�����a�X"��J��d�Xmv��5k�%�ߐ���e���;����=p���#GO�>SPXT|�ܵ�%7J��+nޯ�yP�����M/�[Z_�����sǗ��:�����W��7���WN\\�]\��4�����e�TȠ1h���0��0������!~0ևq1q�����7N��+�ߙ��%���Uf�$���� Ý�&��� и,���aٓ?�����z�8�K>�����S�,���x���]K3?���0��ئ���nc綾lJ�E�,:y���@D���#�n�F3�{�O�y�z8�R|ru*��
����;�+4�뻬K@}��zx����.�ν��l<Z_6�5�B�quJNg������T��w#��n���e|WB{\����S:w�p�ݮ��9����#��zs6~�ŭ*i���k�*���g��۩�!�u�
t/��.����]D��jX������Qa?_�#��n�Ko�eG��W�OO8�#�v�:�ڵ�y��}��M]�5/�ugIV�ʊ;&����m�pC��p���̮Y>j痧��#��.�ÎE�S��\Q�]wpl�?~t?k�����9w�*[]]B׮��cq,����"<#�8��F�l�����dCR���!~��n{�1��oqy���1���[��]�`��L���%ً��E=�@>�qþ����I3��~���j[P��|��pK|�����|vU��ٻ��9���v���� aNAР7�c���3���Y��'�kj��R}C�7�����)�6��V��c��YTo�x�<#\R �f�z�a|�;�E�{m`F�KۆΉ�n���v�?������dw��hm����*ã^��4�{��_�bE4�� �����тs۶~F���� Rg���.�mԣv�Y�͂u������S8��I�^:e�µi{�8����g��M�����	�^�AP���7;�{�ى�m�;����pq�����#ƀu����xY�4_�lF����j:z��H� ���Q�L���m�U~$�D9����c37�{��O������v|���]+D*����yE~IJ�w���mV��s7��{�WU�j��4�ܱ:e)�1�������?�?r�za����§�!Q]���7(�^z�Mp����&��p(FRz	|��ur����̷�� � �l㝸�L�:�����CoDV|;�=3|ݬ���'�m�-[���G���u.��u�(�o[vS�.�n�<a�����3�7��_/�`9}����G=�K�&C�$M+�-+��������s]E�E�N����;��D����9H��;��b��k)��>��҄Vo��QCv~�ta�z}ޞ�.Ͻ��¼�(��	7�)�K}�p�sBe����'�c��R�䱛���3e�V4��K�@�����7�E(�*Y/�8���3zn��Qߎ{�fwx&(�)O ��ޱ��w�5�Ӣ�x䡅����;��5�v�ߵ�m/�Z�#;�ܻ�`_�cem��-;��/r�|��yg�l�ur�'�n�?9|��jPPR��K&��o�p.DX�v����<���R�<��z��; I���颱-�6��ζ��Lᘈa%��/SKҟ-�|Y5hͼ���wҜIj�=;t-s݋A���\��Y�<S�yᴯ�SWϫ�':�/n.�hJ�3�Sk��a/�~���n�o'�^��NZ;�P�Z�t��������t:�JD��kkH|�h�x�夺����!�`c�q�|י[�����*���vR�R���M���,�}kL�C�\lu�Θ�ծ.��^��uh��I_2f��{��^,���)<�:ލz��٫wt��g��֚﫩�&��H>�9����j������l��>�|����͐�.����,O��H�p�ㆴ� j��_ꮌ��<ô�e3��W�9������zg���dp�=z�I�%��D�v?ak��u�O�GD�a�v"���	L�@���#q�y�9giR��jV���s���3����¢ȓ?�^t���$�v<�T��h�|���S�W����!KjA܆����,��݁���ON�~���#O�9�D�W�膝�pO�mMNq��Xp1a�nD�ڬY�G��K���4�o��+RY�^e���~����;���?R��#}$�%+b�S6�'(�Z��:6�.�i$����p��n�݁���o�J?P/`O��1!=��"x��FT;Щ���G��dL�����z/�����r?fuu�_{gE���ߣ�wf��MO��h�y0�>tQpc
ص�7)5u�$�Q��u����-�*��m���+_����������0���"}������~��3?uu1�����͟T��w�.*4���i�l�3�X�j[O9�-	���>p�g�Á��D_,>�dIk��gm���Aƺ��s���
�WT�W��<F��R���|�u�˂�G%����[/��p ��
j�]H���1�b�#R�(~�p���Y�J7O
�X������@��	3b�⦦��m7�'dKX��hu��W�ꛞ�^b�&�[s��oċ�o9��<X�`)ö́9��"cKBc��M�6���K��w�|�]hy�=�i�:���o� ��XO��$���k����n	���RF�Q,^(l�S`��2�q�~䨢+�~p>l��7e��+�Pӊ����Y�;V��1-���2`������@i���&��l[��g�a�s��e�KZVX4�M>Qzיh�3�V�/�Ԭ����$J^����K��B����m�l�*����I�Y�gLi[ٴ���Ή�]�e�ꛗV30�-���7Ī�~pW��	p���o�3���;���o'L;�Yok �$�
�(�="0_�[���8_p=n?�e��{�QK���%�����ڼ<�u�t��>M�Kz�>VP~qe���tZ��R@?�Y���`���hiN����\�)IK���soI��s�<ٶ�Ԃ��ߢ��r:N)����-?��U��ZҲq�M�bRؖ�w'�z>���p�E���y喔����!��[��[rVo׵�9z�����C�.U��z�bJ�TB��A��U��e��UM��ݙ���ĎSn%{S\�\'gi���E0T�tzĹpTḫU-�#��Phr0�׊��Wyd�xj��3s׶�[���֋�G���E�M�晼����0�z�}���m}����-~�/��w�ܹ4p�B��o~�3qc*��c�֔�����w���{�=D��fO?4�*-؅;���+�{$�zn`�� �	������W�$N�L����=�E�O�^H�5��ޜ����f��!-�V=-�B���W�I(��ll\NO-�xj�B[��ӄ�C�������pl�K��\Ƕ]��c鵓c��1�i#�C���
�����i��!s���y����)gN��*�8��ǜ{�����³KN�o�Y����޾/a���/�S���w1	s�nu8)���d�]c�.��I�Ԅ�a������q7^���u�1g�%N�l�N]q��`�W��Ū1����7Mώ�[��C�1̜@���\i���s���Sv|9�N{��~A�nk��ޘ�mz�}�4�q�)� |_��/��T����y���nC]3�ٲ�'�]p��K���ۙ�H8 �K[:皧��)�ϓBW���`�R?��z��z����i$Q��12s���J6{�I��Ŀ���O(Z�@s|N\��X-?n����e᪇��\���\~niM��6�����)���(�	��4�ИQ�s�[Att�ضݲt��ǀ���o��h��O^x��f/�5c��S�c��脛�ao�>���^�0�Cx�2�q��Ud�� �Ϧ�[Ʀ��Eg�&+'�J�]��wL�o�O�xj1iM�W®R���vɤ��.l;x}ăbEs|𬃃�_綜
%}�u�ºd�|X+����dK���d���M˹�n���rl�y���o�y��������)w�o��k'�����tߚCXTS�<�P��gG:s~��#����>�[/`���o�=}�k�~�/f��Hk����f����mN�}:�'yl�E��q7Z\�WJR��=�T�y�;�w� U�~$g���hK�����绾� N�wŶ��6d�����bG�ڲ���%�n�ض�ɧJ�:�PwGE=<�W�ݹ�*�v�r�ة ��|�>�ZvƘ$ɰ,3��c�M�y�nǠ]d+w
Z�9�X?����yފ|�5wUDӖ���t�8�+M]��N`�(�~|9A<����ȫY�e(��\�|���3-�.�^�4�H�� ����ˮ�� �,1�3���L\���~m��?O��xQ��=���Ta�}��Dy����H���%�ʨ]���6S��M��t�=>tΪ�)���'~������<���/W;R�y6��䪪�x�c��O�lc'�Ď[�ea^����[wra۞Mi�ILH��u��QWH6M%.���?Jwm��V�ϋ�^����߾�1���o�ظn0��Ƈ�}�>��Fo��<uq�/c���ҍ��7�ig�������_��}H�uߵ��E�˦�:�uI�5�p xR׍��xe}��\��,�$EQ��P�E��|�::SM���/�mO��;z����s��k��Xn%�%�x�>6��i��c����َ�h��M�򡸑N?�v+{T�����;Γ��-��������Ku��y�ĻA/���Y,�V,~��t�����;#�＆х5�(eC������[逿pyqL}X����_��q
;^0 jj|�x��������=3Ù���+�ߒ.�[�sz��hTF��WkZV[l�"���>�N�ʌ�=�N�����>@2� >f��3��������7��=�MmI��M���@+�|��ޭH7g(o�t�tX��,�U�)����wᓒ˳�3�{���G��$xYĝ��h�{Y�����6d���%��ʠsk���$�V|�VJ,�w/�l�M����h�	͗��ީ��\8�t2r�i�Og�[3��GÝ�+&����'H^[2ߏq�r�=�W�=C?InK��kKi�O�����6`lv˪��R��0�"�b�իǏ]���qJo<�)�+p~#��I[��Ԍ�̾��qh��L�����ˋ�$_1���Խ�X/`!���܃�'#�w���u��{/K��7�?��#5cJH<UN>gd	�{��fGq���g���ž�qz{�i���#�:��c�1ߕ��v�n������*��(�^�X6���]�b�'Ƶs�룧=:�i���M�v��|�d퉪�)#.�n�Z�x����ũ�Y&�KZ���嚳 ��37	`_��wN��)γ���W�ߪ�q�N���֖��Fq�ί��aA�!�ǆ��,��s��1�d~A�=N�����*��oyX�u��I�<�e�.(�Z�ٲq�k�=�$��e������!�����~ �X�3؃���r���{�o�c����o灒��秏m2�h��#C�nF�����Q}��˺�N��\`��B��_4�/���9m2�QS�;�)k�_1�؞�oÄ��#����u�i���C��E�WϦ����#��\\wx�7[����Z{c+��ڲn�N0�}%}+���t�y��!�
���O�tKd}�༴t�ܙ*Kyjp��#?�򽙝?;9�����z��X^�������P���H*^1���+*��z�%HU��5� `��PT�Ԝ��>`pG��S�a���BJ�O����|��ڃu�V��J� 8-��.0��>b� �+�N��l߃�/,*�򘟤�uI����#N���V^
��܅��G�����k�]c��O�O�*���r�:�s_����U�^]������&�w�}�}�Gi����#[��. ���\��K����o�=�𨎜{���>o���_���w7��P����M^���f~��h���ܹkdސے1w�Wʚ���VrU���N]����Xv�и���pkPS��L:��~�|�RXݓ'�.��mlI8p�Zv�x�����[���'o
�X�tX�nR)�'@��Q��n}��-��G��/f߅���];�DM�x�f���#?�̆շ�{��T��Xc�����!W�:�Z'Q"c�RM,k	J�RMW�-�"�앃��w�ؗ������mI��e��{����.9��?�H�1u"�a����i�8C)�ף��n^So�߷��z0��r�ww3�j����Ɛ.�}��t�!"{?O�2I'��K#���;��{�/ݝW�T7a�s�.?��,����ځ��y<h���;��H���V�r�|�����g6�,�]�w���o���WS�l>y�\�c�]�TS��6��=��8a�&��YaļEy{>�fϼ���s��?�����3DQ�zXP6}�KF���폰1���C�ϾYp;D��Zr/�J������K�q+Z��y�q�������:o"�}%�7�t�ї;�&`�'ѴOe#.TLr[�(���%�u��?��x�4&x,���T0�w�H��}��0���Gb�N߭�~��C�w�q�)�2tkx���;���\�/��t��A�O��:Q���PZ��H6��h��ͥx4��a�Iӥp�	5�+�MG�z���=u���ݯ;R�8�a��>=���s��-�>6 ���
��-ś�l�Ư�;��x����s�l�]}�k"��VD�U������[�6{�@�_~��^�O�0?�[���R�`-X0k�4���k��7+WuDD�h����f�A����MoH�Wrm�w��o|y���r�y�c��?��.��`���$���U X'7]pǦOgoo:4� ���?�5����i��1'�F�R'ʛ�;�j!��cn���C��Z9�v6��G]�sp�p��02�m~�s۵�U�Ƀ���ܽ��eF�btɂ��;�ﱙ���3�Q�����AN��q{�������w�y�SP��G|�0�=����8�&1mp�Ɋ)5B�p䷚/�;��+���	͸�7�O^�1'4��=�u�P ���n�wM����@��|�W�v�=��0w�\�}-}V}��c����b�I�cV����#�Y'��L���JwZ=���nG�e����/�`�m-M�d����m�+��p���{8m8W�}��h�����a�-[�y�sq���E.���Qx�)RB��H�	|�3e1ሒ��P�-�-k��J	�=M���s`k�
ZOױ��^�Tꐉ�����jB�>̟0l��{~ݣ;N��{�쐉�1�n{c��!�撒5ύ�kOd%!�Tm%-��u�KH��7���B<��~d7�Z��or睔ǩ�ŭ���vT�Ⱥ��<��"��t	��g%>�;3!ű"&�Z�����K���[����.-�A�,�t�#��@�� ��פ1ao��SO^�%�<�.��^7�ʭ��������V��^��=���׻�����j�G
�C�
%����B�>L_������,�n�Uzd��B�͝�nv�z}I�a������S�F�=|�����^��zL�3ZV�]��ɺ�W<�'\�m��a��4�:d��H����M��oo�v��k�܋��m_�}�Okgq�w^I�WD��sx?����F�5`��SR����jŉʥ��n����JY��O��{О�Y᯼�y����X:��x(0DOy~º9��E�e���X5Uj�{Ҷ��^i5�L����b�t0������������/�ݮ#���[�s��.���ʌI)���w�ܫ�>�&�Λ�����"p�5	���E������#��F���(�n_pL�\���Fd�F����=3���Lk��*�����b���4�X��]�k��şF՞{��ß���%M|��G��s��C�<k�6>[��]�Kv��`.tု�g3n��[�bY���M�wi�1 F�r}��{��s���[۪?���׭'=�Nd�'n���ae���Y�kuM���BJ�mM~����{�Љ�Q;���0�]i�@~;6a�[M��Բ���S��r�`��e���^�5��y��o�~B\�e*��4��F�-@UVL\r-c��k�)<�}�	����o��iESs���)qH��*�ƍ�fl��	��7�*�~����!�+oh���O�z�[ᑪ�O��K���*�/;ud�Ɯ��Re�Zɔ8��th�x�ΐ���A�0͑-��6?þ�%�g���RU��������c|2�?����` .s��A�_+%3�p��ݨi��P�ዿM��~�j�Y������Q�Î�9�I��>���䐩��b�ȝ��
���P�I��I�?w�^�^��#�����3O����p��`�X���/?��#��N��9/W�L�:иiO��S�O�m�]�<����Q� �?�J�^�B����-.����Z={��'s�Nu���~vUɦ�y�X8���*��{���;*�yDpcc��E�`lO�~rq��XP03k�g�c��kn@,９��.C��&�g�-��x��'�Y�Fզh�Y�h�^�j����q�zݢְ5�s���#�F�^�P�V���z�s[�z[z��-��_-?�\�������Ϧ5IO>��TS��I����+W������Y��d8�����C�W\�*='� ���Q^?���2s͚��2���$��3��X����cf��2~K�ӄ!��ŵ�vF��X�b-����%��}̮`�����������*l�3У��u�[!k�:��Ǐ���+'��N���r䮾��m���4�'�q���9��Ys`y|)JFL�[��,�$�\�������k(q����2\kdW&��9�S�Z���s
�9�CNKH!V�ˮ���P�_p2]�}�����w�e;V�sV/`I���X-�R���l��цO�|D����Ek�\N ���o,su~�f@�vot�ҫY>�+��^mݞqJ�8���[���A�H����k�n\�e{U�DLz'^~y[w�Ρ��"=����'����G��v��ѯ�i���y,��F��Fȯׅ5���s�\���~~
�ʊ	�̻�j4.kg�ߔ�[���˘Zx���S%����)�=��k��7����+���mY���|ܷ5<�Pu��3s��o+�ܢ18��H��J������q/*�t�;�xqޙ�ƪ��Y.E5ک�,����Rm���S�<�q@x���6_y
�Đ�:��Z�p�znם�]V����ot�q�6��ۮ})Fd���zy%��^<���~O��l�͙3��?p����i�'��c��M	�'��<�&��1	�OrK=�f�A��=�U\�Q���i��qCe~HRI����7OQԷ���̪gx���H�d�<M?Ȑ�c_��%�aP/`4<�x�p"Udx�p�k������Ϫ�M�?n|�r)����w�n; ��?�{Fuh��ߌ8,�cS��n��+0�;�Ƿ�f*�t'vݿ�U�>��Ҏ��mMMo�[�����Mł�×�/�<� ���������)�u�v�,��Ͷ�|��L��ȑm��?}ų������L1%���ouF-^C���i�~ptQ銍����sJ�'��~Vwq4Ȟ�����t��[�<ؔ3���]�3�>�-a��FwՊG�.��I)K:�<��i"{���J�[�g��:��k�kW޲_�;K~*}Vw�c���D�G��3����-|��-����r�	��χW�*��Yv"D��6�[4��*�(�})��\�֘�o������]X�w�h���!�-��垕:���E����1t9�;��J|�p��m���?�9�)�\��
[W�}�饼�E��e��~U/��:���������m��VF/ r7�d�����-{%OLےr~	�W}g�q��<M�]�������t�np���p�޽sz��6�(�v�LV��2V?I�;gw��|�[��YU��!�0�P�_�=�{��-�wm=�:�2P�F�wD�]�\�e�d�{tqi�`a�sm��.ע�ƞ-W��/dt�,�L��U��(��}���Yo��86|U���%0�ﴋ�L�%c�"�W��h[�q^�z� #;mrރ��'��?&�RN �9���`�=�v�[.�r!���F��h8��"i^h&���A�SӶl>!sNh�:�nV,��#b��	�7��$ο8��.t~�jӾ����� _��|���ǔ�=�����eo9�����<uܚN���"p�gZb�A���q�6]�y����3��*�Z�O���Lb�T���􃛪bo}���sq���i~ɰmw�:{a���,��s��v�ǵ��^��v��N\`m;XWyx��w��y,�JX��4.�v���HJ��y*|䊶���m�:+�e�G�4�L��dԖn�*˰��kY�3��RL?6��H?��H�Ln���<�.2xU8y�����w|�x=-r.p�fyq�!��<�c�ꖴ��$��7e�>g
Nw-@�|�z6�}���m�.Ys�2���K�ϼth߂�5E5�x_�ˌGC;���	�5�e�G��r��d¦��])�)�gM�8~�̢�- ��̞�X�Rw�e֔����Ӗ^�T�	З|�W����r����zyߒ���  �5�~���K�е�-��7��iإӋ�^(J▊�#w<ϊv~'�"+�Q4����s�Iu�qN��+^�s�a�^͹�d��i���v/{@0�k���6��1|��Ob��Yӆ���|bLN(]:������5��Oy�>�3��Y�?ݭ��~0������A58ΔU�Q)�'��G��-ӈ�@���&�8v&�G¯�xc�n_���[�B���5!-���ܯ*�ŅLև�-���O��O�����/�G��k�6�Ȼg��_��№�k�n�}���m���؈-�����u�+;���_��\���]:���^������m��1�̌8O���)����V㏢���KyFϸ��9�F��Q���>��=�eS�OG������$���k2���şv��.��W&_z n�l�w|νֳ�����N�K�6͒9���YЏ�P���J�a���j��x��N���11'�!6?���ˬ��KZqY�F��t'��A�_���	>��6�ۺ���s?t�����;*�,�#`!ѵ�֢G�ŧN�N�I���᷶����z���R�p�d�3�wg;�o,������;A?�{�Yˮ5����]f�y�7��^@I�{T��hTnP�%�{�zX�F �Uu����'��4���>Njr�!�]�i����OS�Y����&�v9N���ҵ��_�c���T�|0������w�{~��L߸v�2H-��m�����n��pZ�$�z��ǯC���}�
���焿?�x�&P;q��o�=����,��|=�몸vYHc~��`[�������:k�Z�69:��>�m�t+L&}0�5�It1ҹb�d�A��` �l��5R��Ǧ���ma��݂��j���o�:��넏���������"@%�a��F'�����z�;
����j�ε����� 
��� (4��#�hךD� ���wv���qJ�I����:��̦0_߿c���:�����kj=H�w�W��EF��$�J�����|ap<�£`��"�G�Q��@��������?`�kP}���G�IE&]G����?�{7��6�7!�U�7�}���}���|��~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~��5��Eb���#�J�fXg���m���m����aT� ���v ��߯�J���^��t���������"�����_�����/�{H��6fo���&@���]�B�_���q��{O�8���Z��<�@��Rq*^"�a�Dvv�^A��とf5�d3!�1���B�`P 9�D�"M �M��Q����`x�Rna��VKkaƑD�F�"b�*�A�5��QJ>�d�G�,�J���XȂ��Q�
b��,�"�4Qt$Z�QY�B3KıxF:Q�G�đql�\��bHt�	d�Дz����D�X�Ç@�y1LGdl���1�x(��#�������k�J`����DA �o�km��&�T���qLt����xD"$�ҴF�aIb��d��m�X��E�
b�Ej6�f!BY��%)mb���(#5f�.e�cQ�5�n�P�
o'��xV`�"�(�B���"T;Vt@8��D��RF�IA��`��	���ʌ1��h
�%�¨&�F.�Z�v,O��$(1JdW����Pi� ����∃��ydd$eb��
d0��r���$���H�����P
���[h|
Hd��"`l��+י��a$�ˑFZ�f���3� T�����|!VkG�Dj�G�a��L�ԋ�j�)���j�a�f�D���V��
c[D	�KB1�j1���3y$C�4��P�� �(R�D=�a�D�٘��&N5Q�t&W���D,����`H�H�!qL\,)�ȦID	�j3 ��J"��:FF�,�A��T&6.F��r�`��FТ�+4� �K�}7�)!�t��&��Y��XP�D@	R��JE��f�]"���%@��*�Ђ�h�F���0�4���<��o"��(	� �F�E� gB��jB���D�U+gRXZ! �"�24W���x�I�4��MR����B����p٢�`t�� f9�rX��E�Q;�ĳ-d��'R��r�<*H�У�p���3��
F�]�5GE�"�|�Z#W�PuD�Ȓ���@�>.P�Uۥ`�.��7�@5�����8��&#p5 ޤ�9�6u:V�@�yD1g��1=0FD�Ea�<��D��
�L+H&@G,D6��5R�j%�
��5R+�C8HD�Q�p����!��!�*
QL��bY�2��cř��B��DE�l�چ5qd$�CB"a���Uh��&Ή2�x��)�;M��#��Y��sM|M�&��$1�
ˆ��R�Eņ��1R��b����b�c�,Ԇ&�|������D;�)P[�BF)��f�L��F�QJ�XƃJ�b4�$F6�T��E��6�+�9�
*P���2��q0,y,ΌFPIR,4!1�
6ɦ�),��3���m&SI�aC%b��h��(�h(��cX%���wo��̾Ǖ4���!`��'C�� �K 1b,�e�lR���Q`��z�����
���"�ݵJ
�j��"G��4�YT#FP1�$�؂ֲAX�>Ȥe�a$�� aplߪ	!r�P��S8`�N�T���H5���J"YnR*(���i⬢ ���T��\8��S"uQv)u��$L�C�PP�����@�X��xZ�c���h�D(�[���(6�$e�H%'B����rXd�%)Y�@8�P�H]k@j�j���RQ�X����q4�P�b��HG�35F�Jf7�l<��#Qp�2[
���@e����R�����(&�ȵ�c�l*͡�A6^G@�-��D$��s*�����F���b��H�j��N"T`X|���S��T<�ͥX�b*N�[q���YNB�ih�8�(�W�j����A#�VpC��Pl�Cb6�a���p��6��#V �j%l+$�ቹ��� ��v�G��j0Zʖ�cIAR.��`��j��gƠdl2M�A$�H7cP���lS��u@��G"�t�l����Q�R�5�ff�l����l-��E�aD;��D�(�O��U|����l��t��G�@#�-��if$Mc����,9-
�Us�PD�0�2�CBG�l��'Z$j8)'��:��G�%V����Ȍ\S��(q������+�����6YgP+)@""
#0�@J0�ȓ�h��Ad+�B�o]��c,P�L��j�����c���4c�8-O��1j�Őit�ȁ��2Y\�����"����[5� �'�J�R��Ǩ�4
��w��)�V1��2�M�$=L����$�u�I[Q8����@j���t.���*�	�&dJ�&�j�t�IŲʕ@3;�ǳ��(zD�Y�78�$�ͪWb1�\7NȢ��P1����",���Q�X�L#@��&B�@(�X
�e�Fq�A8�	Aj�4#Xb@R�R��j"���b��r��"�T�N�)1@8��s�:=\�X-(*�Kǩ	��C����8�R��h���H���)�@	��	 V��3b�(��ґ�f�*��"I��(H�PF8�(���j|�HnG����	$���@=�G����n�K��JXp�Y�$��tL���:��l���P����L��bS�5h<��(�x8W��ڸZ��R0�� �Y�d
Xcd�H6-=P�\GB�٤HM �Ш�|��% $Z)Tl���(nV*t������� �����q�:&-�[2+�p��Io5	D8b,�"�bu��E��}jTBժ�~P ƇI�F��%��QDzV���rr����I�B	ȀB�  ]�1��L��a!C��	�T%\9$�[�JNoT��0^H�h��� �j�������B������f�n0�M,�Zk�ӣ�(2��F���H�尢�x+�C"��.�"�7�Q:dL��G�D�`��@`*�&�2�����	|>EA�d�J�u�%\�Nn`�hl�Cڢ�80 2#��j.W����q\�L�)U2m�g���(���I
:=���
!�g7�5:Q��[�[ D���L�Ǎ�ɀx����3�
�8��>
(��0"�`����pF�E���@�RG�G�y� ��ǒ�PAH���A�0M05C���pZ.�	�D}�a�3�`B��5���I�Ehv�^�`�1M� e��8>�e��0P�\���T��!�b�v�D��)
��&��Q�#�E��X��f���6�'�`�b�
^OFp�|R�L��+�6��L2����J���'��\���I�q@�̡�q�R�$"��2Łht��ų���`NS"��qz��$�������F����BC�����
�I�R��X	ʄ�uK+SA�&��`�mr'���IX�
I���ih9J�63Y0]ʓ�-(� ������v:F���88�� Qi�P�Mk�+������"�Aj�َ��X+1EU��(Hg�*�T��j#aE�H��@�q12]TiV���R��8[ˍ�iuP�le�%VVA����<�#Χ�c�A&����<�H�u������hdT�R�'�qr� �#F��$�J#ԡ�X0�dƣ�l��Z�r(��pt����4��PX��(Ң!������b�Q(��� 6���w��M�8YA�}�읢V�5{y_�ȓ@��j�R8���/��)��;8��_���fW��L�zݾ����iMm��
�>�~��]�[�[��#��-h~�Q%	1��!1t�.��疵�3}x^n!��ל��6&�r#`ҰT��s���� J��c/??"�~��X7�H悥�"{�����~�j$i�#"�+�ZHbR	�T���;k�i6�K�/��ț��-j`h���Wf����j�����xο��`������ڰ�I+N��.�[9�=���4h���>�9�J1�H�H	�Z��9^��e��2���Z4��=�k����lF�����&�AD��x�Ϛ�� �y���6��Jh��ן��R3mʾb1<�;<:,�RB~��
�@R��?	s���v6���,������v��L�"���ԃ���W"�X�6�7���!�qSIш�%XgSXǘԚ'e�8��)���q4�Wۖ�eU�}B�^��Ý|\'�I�Ċn�O_�z#^Fӟ0�ciz���ķ	�p�jD"����-?��Χ6De�*�
��)�~��F*�F�5�v<x�W�y�OW����Bw���{E��2a*���E�VZ�.��bPT?�qS��uXX$�z5�2/W|�κ��8g��+�b�71��f�f{Bdr�~���FОY0����&M��:��tN�M�$a&ay�������=-��/-��R�[_�|�^��wX
4����|sO�)o���h�>Fu�$ո�q��&��� �)��ٮ�\w�t�/Rt��`��N�y*����J.ơ�X�]�U��/I���N�Ά��>(M��}���pA�|��~�;���nb/A��t/$���
�Vy��7�#�����c ƾ�HS{Q#��y��r�.�����u�Zċ�#��$L�E�����q N�ո�."�)��éf48�P�X�@'xK��-�DQ>�)��0c��eV�mH/�Ƌ�D�X&L}�@�m�F�%�瑵��^�^D�7����Dn�l����r�1K���$÷JyO��ٛ*ը]|*�a9fл^�?f�����۶�ꫡ��BD�´)8c~ng��|��r1�������U0�m���IҮN7�?�,��rL��J��Cc��e��ǡ��T}91�?� '��>_��Y��4�,.fD��O��k߅t�l{���!�a�k�@�#2G6����qƆeHVC���8p翽O}����q�<.<ײh���_�Z�,��e���&�� �b���,(v燩�aҨ����"�E�|h,�,��D�t_O�,�#�h__7lH-�BC��C��m���Yt��R���ߴu�|o���r�h��Cq���R*"y���N��M�o��w?��$�||����ޝ(%��Q�[��_N�*����2'���)s�l�ͭj)�rt*�#,���:��B@���S�E����
T�HΠ�s�5j��!�ڐ�t0��C�A����xQ._�I�Yo×����HǺ�nӫ��,��a�zM?�Xs,��[rO�1�J�*� �P�q^)�B�h��=-���%DT�{ሡ��Η��'>�g�G&����ô,���_*ȩ{�u)���Ɓ����5�{�)���\�&�ߗ@ic|nۿ^�Em���pA/?�κ<pϋU��bg2�6���C>��#O��o��������)}�Ӎ�� ��/�,<Q/H���ܒfV��w�V���&���HT�p����23ƤK��L������������ν/�������J6t��*?`��դ`v3	�$a|~iϸ�k�پ8���ll�.�H���f_�E�}�l�V�~"�<׽�:D�������~��R8
�VGbQ��9�!D���I9�&��9�l�r#Ag��D�R��B���ɠl/+�0,���O\�CLuW���x�5������E�s�4�>�?�	H(C�IB+Ү��y �Ƚ�2�7B�L�����.E����*l�����p��0�Xl��c����'�>�{!��=>r�G"�nŵ���[� ���
>�¿��S�:��xV�aq驼r�`�_Bg!��]����Q�?� �q�}��4�}�Ds� �-�b{IV��!X��%�{ɻ�:8�[�8�C�w���N�O���I,[>u���_~�q�G�?j�w��dA�*��0��6���d3R��A1y�Ů�����눬-�g]փ�����^
^�:T�����n*�N;�}}$n�s+G+�*��6,`��K�y��[�+#��J��;_;�5�}@]%�����J����{dݼ�ŧ�'�J̻u�Fo���@Dc�'Z�'��[�轶�&�F�&�CG�?D`TG����d�ޖ�1б�S~`�����o�GW>Ղ
 �D�b��-��,FZ�H�tZ���ǩ׷PR�`(Evѯ�5��ky�N�j4G��;Fp����qhx!�puB�����U��W�~me9���@�=��^/�i u�t[mq9}n��/��z����Y��p�l=��J�B�<ۢ�o�Kn���s�
\������i�_d?�����H瀤dɌQ���B����P��!S���,ą����M�I� F����\��r'�{lS�C�Y�|2O�h%c��(J#6ʥ[*���c�����1�j����GTl{��Y�K�4+V~� ���'{��>�w�6��K��������,&K����X��a(��EI���z7q �o�7�Nu0�Ÿ�V�R�Ga��5kӪ��?vF�`��P?*:�0��X��/4�bB�*�o��Pb:M�I�+���+��ߐ�8��Ø�!J�?��S|��O!C�Xvukc�t��/��Sw�*7�n��S����D�u��60��.��9]��ckD�K_�u��me��7Ы���gZ���r���M(6/��$��}n������U�zd���7H�.K{�lMĶ�]�C0MTJƁ
H�k���l��ҡ��G5z�:��6�5(F���/sʥ�A�s�|SP��s<����~���x�;��̌�3\�t+�@Id�I�gm����D_��#Ά�*z[�sMs�ph�7k0��5�o����=�Au?�~��ռ7�IZ�t:�Q��^`�I�D+�D�:yMɻ��sÖ���  $?6��l�Px!����^r[0�����7���!{CCXk�V�9�T�����~	�iRH�<��&��q�P�{�JL?��Q/�A�����u?D������ɉ��TlS�TUVi��3��y�H#���jq:0�e�}��%/&L�Ǐ����}62��w4�Y<V�3�-rCШ���1� )$$�ؕ�w`p';�}�����G"���o�ئf��G�����:�m��ih��
�,x��P�]�C�	].D>��W�!vH�>�âE8��-��#��{��&'�w�L�#�@�;���Y��ТP\��|�0����̆����[��0��l���V����5	Tb'E?����Csvߙ$huD� w�LA�#{v>nP�8F��'�m�47��p'�r����"�������wJ]l����4��D��:gh�|����LSL�pk@�������a�B��CJX��<t��Z�Zӧ����N�>"r�1_An����{�|���@�vG{��WG���V��vG�gf��ɯC��&f�LHrR�HJ�&m�y����0X� 4��wh�5H�T˺~�W��/��FT�|,�4�1�*X�v�{���P)t,�C�c�k�&[ٺf,�l�,�И�C�?�&L�Ph���6���"���������y̬�-��SЯ}��_ql�����3��ĉ����n!�~@ڥ��Dg�X`���Nbf�Sdi��b���P�#�k��N�B.S���;�v�3���6�o�T�k_��.4��'�,��3+�%]���]�+�W���mh%���}y�9T��0�[�����d��9Fj~���X��
�&�O}O�B�:�T�i�I�9�C*�����jIe�Vo��V�o}Rͽ�N�N���-�\D��[�`��ѳ��oV�>��.NMN9r[ڇ�L,;�m��:��1Ǹ��&��3oG�2f�(�����n�#�fϑ�Ð&�r�����ﾬ8�!v�ƴ�/�,��8^/
��j�}e���5��\�Ζ���Ao�G�1(e�����N����(����{�ٖ`���k^T����S�=.f���,Fe[rA\��։K-�nV�lLQĸ�\�5�__6��x�-�2���;Q�B�|^cS��n����{�=-z�?�	�C�����|!G^�TNmӎ�~}!�){����)4�y�����$U�)���R:b�7ѷ�l�ȓ����3�A��ѭww�U�y #گ�.i��\n��3�]�YP�!���!�R>t��#�N�ࠅX%�+��2�+�ylF��`���zQX�ص@���Q$T֡IN�+¨eCVr���!7�d�8��4{��HmQ(�|�<���sC�-���G�w]d�a�(�[ zi�vQ@���!����7¿��W.&!R�~�";��Y5 ]�o���5�}KV�\�}Ie6ξz�|���Z��Bv���>��κSL_�f�%�A��;�!e&n,�b����ުﹰ�(�s���u�RC���9]X�Qo��7b���Ђ)��o�}�n��<4[c]/B8X�3��u��/��1�w����Ѯ�����6�����������z�44�������N��*T�p�e+��M!�]F#��Rrd3��ҍC��em��?�8ݪ�#�d�̶����8F� Y��vM��w����nBDČHJ����r����Q�G>���~{��*����w�;|�˳�U���+_�ҎzS�Q:嗈�!���%!�"�x7�i�RD$9Q�<�ȧ�3(� ��Qi����?����	g�d���g��c�����(�o�PQUH5	m�v���A}�NT;��b�`Y�#�@�9�gp됅Y��W�$������jS�/����z���%��$נ��fC�O9��N���+�m�m@�����x�]��8�*'�A5X׵�����&�[{�_��E{,ޤ�<��;�jݦ"��`0}�c�U��`F�6:u�MX��өj��}�5���/\`���~ep��Z��2��u��~g�(^3�]�s��/ib�6��K%[$�\D�ov��p�a�jP���	�t�nMW_z���� �~�8�-9(�n��~���n���5Y��>3LRI�Wר����d<�������T*�3|���YV1`��_�k�{�ί�,��S^ۭ������z�聀�0��PE����- i)�{T��`��:���p�˯)������:���<�;�_)Y��Q%�< |e�#]V�ꁠ�+r�o�Į	 	<N��8T��$���¹��[n5τi ���X�zN/ _����o*b�U�[b	3�(��	Ao�Et�u&�)E��T�h�n"���$n3��(�+��_��x@��14tҝ��g�u���2{ |�c�~�c��L��(�9��:ʼ�p_�\���*ywbcRs�6#�=R_�ㄕ�
��ήG_ٌ�%�`BuEe�`�l2Jy� #9E��~�|^��O�(���ū��w-[D��+Q�P%�^2����N�_Pr3�H�K�Po*�D(C1�ʐ�k��3�o���̣�U�f`� 6�{X��0f>ܺtk������)ֳ\:oV��#~������j�f_0F�mH��Fd g'I��N�4�^m4�#sē���{@�/D�>�^�3�+N01_&�8a��s�h���p�K��9ص�c'
4<�[(/�����]��!q,H�i�EA�:D��Wm��|����2<��/�4��Wr��g����Л�_";�#��$C�O�d��~����בX��w,��"���@dpq���i�$ "�,�9�:3ד��r �Tc�)O~c�w��_C�9�m�����K2�|�X�!�B�m��Ɣ��]�+���f�Y��T��31�sL�]s���-�?��}X�|�svXĔA�ǭ�Q%a)�G*������ia��F� ��3�1b��n�-^]����Ö|bQۨ�J��t)iI�����X [��q�&S����}&��',~I���3�y�,��j�њB#ᚆ}�[��Ǹ�M#�T!����u��%�?��2���b9�|���M�m����zu,n�Ʌ�Fy�}w���M�M�m���_z�4W���չ�Fj+5X�$÷��7gҶ�>Hą��;_��lx�L�YZ�s��E���3���&B��(���� Vj���i�s������a3&1I���^�Ø0��)9~��#�b��)[��\/�ߊ�Iq�H ���lN:A;
��m����D �>6�e]���~���2���䥎��
�vt���/
�q�e����R�o�U�}��\R�Ln����(�D���`:[��]��; ��I�I{��q8ӽ��*7���7�W1�U��v}�6�R���6y~sAksɾ��OU�i{T:�N�9�9���P)(y�x#� W���ͼ7o�Qߏx�y�*� p/�$8�G"D�G��pD�ۅ+���_�_��1#C-��\x݁�f��Ni����~:�~'�k���@�7��S
r��m��<肚�ύ��X�Zc����C7��HX���06�	���i;�Z٬S(�U&�-9�6鰥ǁ��qfo�)Bdleb�����}����'�>��2�YA��"�����8�F�$��F���:��\�w�&��9�d!����wx���IX�!�8�ķ	�(싧C�)��	j!&�=�����������c�~��ޫ���� �$�r8�L���wK2Ko1=�!�駷�2Dg^��>IV	.���Xپ�i����BB�+
�������N����ܔ<M|�A/�n��c�aD/6�*��8������9_���I�Q���-��� �������9x�7l��>Ws!
�񬾒�1U�~�����j*t�5�� �ZD��g���L�Y�7��H͛�x6J��Q�c�~�q���ԎpkyQzm5�F�P���>J��NpR�
g:���!!uݛ1Z���{����t���f#�oiu�T�QV��B�8�~ݰ��^F{J��\�g:�\*��Z�~���Ք�A�����n��%�!L>�|ʏ�zޯ��&�=����xh|��}��ϩ���.n�Uv
�1�q
Ƀ.��]�F�j^C֙Ĝu�-��o�M(,8���Q৭�kˈ���.�PM=�ǧ��"��F5�t�$�
^R=R��_�́�sAp���|�)Sӵ�ׯ��l�h��@�׳�i@��\)��"d��\m���TWo���5����E`�6��y'O�0����B�&ֿ��Hc�6�z;��feB�x���G��p�SM�4;Bl:�[��5�F��C�݊�Y���w���n��������=����o��/�Z�@�7���Al*��	}���ߠ�2Z4ǀ���a�R�˹w���n�h����sO�K>Idb�#3��3�#!?v9To�u���M�JY���r�Ћ%�.J�s�t��><b_�}'���I)�O橳��+5�J��Âs�?�FyzS~�E�r�g`;���a:���+�:l\.;Hi�B���?S��/��{�{g*�:�C���z�E�9�םy��>=;�K�]ra�M�:0�9&*�e�X���t�[a|��=URz�on;i�1q��Kj�5;��[�g����%�������.N"�;����L��^�JB(��7��c)�ZH#| �Qe��:��4?�o^o� �:�v��XCr(�f�U74�I��DÚ��+_�0$�H�� �u��M��������ke� ��h;IF�����X���X��G����F��wJC���*�&��0�6��`�A�6mS����γ%z�od�h��>� �c�ź�z}6x��� M��%�>%Rl&'�ǜ��8�@d	�]F��Ls��r
 �.}�E�}o}\�w`�T��-�8�Ge�n�=�b���ׯ.E��Ӊ�������#J;�^�)���M�*��*�>65*̓��?P�:�)0`�p�C�_A���nZ_�����ꞝ_���R�
��E6M��^]X�4�Pa��Dcv��6��P��a5 �&G���â ([�P�-���� �E���:<*W��:���G�$�
9\�A��.#���l��s���l�U�L��|���[�`�]-��ԛG��+���VH�݁1x����2q�ì�NLB�OrȂ�9v;���0�;�◳0R��ܧ�7�byKdf����sZ��� ��5����t�{k�����J[�7��EY0��%�9����W�������p_4P��{m������8���1^�%u�hU�rw̟��`dBh�X���"{d�5��%�I͉�(��B�����Q͞��x��k�D�Mܟ0��;�B_��Y��ƭ?<N�'V��7�sͅs����&�!�;e0�
%x�	X�r�(k����J=��Y;؇�Y����P5!&w�k�ݓ����s��g�����]�j�/�|a\
�=5���̠�H��>W9ʗ>��R�"��� B?k)�Ta5)���ӰPd�Y��"-��3�ǂU���@�ԟa�G#��:����0�NG����ޫ�)�Dƣg����^Dw�;���Xz�Q�u����
��X髜|4v�oI��dt㓦^��6@�h.a��p�Zo�����$�Iw�k߈�&�3���q_�;�Ϙt�:\
��z�q��bN���� ��5[	X$�8,�W�6��-5�![H�=��E���`kP-��Ft�j.(x���ܡE�v�3f��ߝ-�AK����3s��S�*��t<��R�{maRT��˯`P ����������P�:K��`��{;�k�[��<�`.c�Es�\�b��.��l�Щ����h�R����s�"�����%gҔ�c���������{1�&-�Q�Ҍ~���s1(������q��|�"�ѦT}	�Z� ��,󏄍'";��p}#���(R	��ڞ�����^�:����\�߱2	\\ǫ�$���Du��#�99ԝ����.�GS���)N��xeb�y�Ը��W\�6��p��U�fKh-�&RQv]r3�s�d�T��!@]74o�qͩ��DU/#��v�%�!x�C�{�^Mx=hW�Q�P�QX�$Hj-��؆�}�O��"\g[M�5���h���9���{D<�R��߱$;[�Wg�Y��O��ٕ�t<�����$W�[�,������h�v� ����΢�N����~���G��K+��A�6�(T�LHBs%��[�
��' �Ϩdn^���18���z;ó�Ų݉��Zew�1Zk˭�Gri����v��!�I\�x^R�)k��r��j��Z�ʈ�z϶��
R��''&�X���l���K"ə&l�v�2KY�WO����ra:��	o���.�<�uJ��1nH�W$�u�P���
^�0�W1����$��A�|��m]�%�A�@L�2.����xxZs�{ກW���Җ�̯�8���C{�,c��~�P���	��g�8Sr�����?�{�C��'phBp妊��H��˞dt�EI�K֡�jK��ߵB��ۆL��]#��y�g7�f�����t��]�d�S�pƑ=�ښ�Wol�	h<��.P֘��*��[y}��!3�b��tͮ�4wh��F��*邰%�Ӓ]"�[Tn`g�5v橻�s�]|�L|�*Ȝ��egF�Aܻ^�7�X�<�ܔ3x7�!�0�j"-�'�SrPێ4uLK�b�*|Ĕ�Β�?ڲ#�v�bF�!��A�+{Y(��/��8���]%D���$୷�zNx��S	u�����oA>��/;�~t��v.oD
�mA��5@��w%J����k�T��&��0��QE��Dk�v� Y`���*�c��=���k�ˢ����Wj�n[w��o����yD�U�/(#��I�!A�H�i�u�9e2��������ˋo�)RT�`|��M�w���a��m,�����wK���������ꭨ�p�"�x����ض�4�FaP�ꧏøI�CQ��N[����3�#�+}���}��M��	�6Y�9���A��.&`]����h�r�ʍ��>j�(��dkc�ZX���i��[�'����t�&y��f��Yl�H�_��Gǩ��T��+���Zk���1�HX��v �]������m������B�tmn�ʦ�*ܼ��qt��df6����t�z+���.�[Hdo��������	���SM���M�Ï��ⳟ��kȿF3_�6���g�X�|�>?siN���f��!���E�@UC�c�Զ�$ ��Rm���F�X�/�.W�ښ@N������/�$r�$Kh��F�t��w�s�(��S���b6����Z���"*�&KU�r�c,!���8Zd�3d2V#P�}�F&�1�y9m+@�s$k�5��baxџՒ�9�i�Cx5�"��H�W' }e��aT��8��j.�o��~n�~���|�f��WD��`���W���z�	���u4�"׽�"*�x���A"o'��` �6��C�O�ک���:����>��d�Q��ݵ`�eJ��4<���F�}>j��K�ٝݺ�ⓜ:ړ�����9�;�}Ow��X�؀r�5v�&б )J,�ɟj�z�T7�������XdԦ"?$�Èuq��#�Yya`>L~�"+�|�}��L�p�.����rl/-���3���zU�!��b��Ţ�����A�R��=�^^����Qgz����@��dP�c�u�M�0bi��o�3ʲ_�R�s��P��.�ӝu��ܙ~�D�\���6�j;y^mn���!x�`��n������#u\�������#H
J=���7sr�Ќ������J��oBN2�S��n�����S�,��,���)��I�ݤ�~��c�}7�>)ߒ��*����S%E\����6�Ǯb���w�qf%������Y�{~�9̀k�Σ���v���`���R�ɠ;>�?'�]%LJu�d_f�XX��RI�>�=��Qe/2�-䜇sT
��F*�� y���Ɉ#,*������-@gx[�����a'V��� ��Q���[�'΋ְ�R���1���k��t�M�e0{�5������k)B�ӆ��t`��|N�������xz[��&`&�x��L���F��'�d9��.�[F
��5�N4ϖ��9F`0���cS�+(?�u�r�"�L��(�nw:��jS��O.O��6�xop0�hc ��c�'��Ҷ���S����q1��!�H��3�lP��M@W���ܜ��M}�S�O�:�z��d�������i4�sև� ��v����7�����h�c)��=�)�s"�`���2��U쾝&Ft�,2�Ġ����'��iT�Z�f��n�}��X�T�I� <U�_�d*JN�tV�oQ�`�{�~M*$u�G��F��Q�TU� �`���BZ���v��i�A�F��Q�n2�#Z���T:> ��Ӏ�"�߬Z�z`���n4��\����s�u�b��?r����҆��Fj��'�;�23"B� 1?���cV�O�͖8�#A����l���a�]�K�_ǩd"���<ަKfn�_��	������5���4Z��d�~WVT�^k��um��6�?u�M��E��]՜=;k�ID.�o&ΩY�}I�R�@���}9�g?�c\S�V)k��m�����5`��� hf�Z��5��qPX-0?�P��ޜ3��y��lO;��>�,��^U�8i
��H*�|� �����%�-��0U<a��=�y��J�+^�k�y�%O��\�g��1�-2�h��b�ޓK\���J��{Qn3v���y�����a�{<�p�#�l�v��+��m&d�~x$h���в�l,�c��P�R�/����q�w�mrz���2Wh�@g�f��2
�Z��:X��AaX�V��AطÿG'-�F&Ջ�pu^���~�Ԅ���кļ��@f���7x��p�w�-���� ��Q�%{���=�(A�U�P��R�,�p���q� �/��Kh�F�
M>�k��E� ʤ�m���<ɟ�u�ȳ�T�	5qTTGc��h���!��Լ���NШը�y(Ye���:-��'�
��e��^̉�������s�R���>���Ԛ��{p��g���L�' �B����7�1�j�+���j�Jꩶ2������<�#�����t���vS�7n�$�l~����m�W�`9�l�	:�}��hhL�A��x��Ʌ��\J����M�'�k Ev����B�!���O��λ���kF`��(г�p]D�J��%�̳P~�/~�݄p�L�{�����r��X��09gv�3�f9~ol$uW�7H����y'�Wc��|�F,��)�0��TO����+��j?��	}s���?�6��9��j�'ۭ�=�N��^­?�m3����i���7���z3~��Jn_:c��Ȣ�hI�y}0�ը-��m~�u3�ݷ����Qq��7A�zcDH0�.��Q�?�*O�+�&��^'�]^3���d� [���O�{X��՜b�ͺ�{��䯼��WF�Q"$b�� �=|��-�h{�k�dJ1�x��v��+����E�U�Xr��P��8܃!��wg�������&�Kgç����F
`|��� �=�8��A�4N�	���,3�4�^��<eN���c|R����$��%e[��7X^=�����*Q;[�(��Px^,��?"�
�� 5�h/��h���o�2�<���ſ��a��mQS��M�8�I�!�K=�F�B�O ����ԖMf����Gt�0����%�n��=+n"��^�K9o�!iW��Wv=9�`�7�̆���3w���FW3�Vs��TZ+=�ĻJ��l�z����,�RX��	~�7>�e�t�Z�.�a$B6��Ƀg�N�WD�����]\��.r����K^;9�����.�Θ+�k���tE�&������i��ܾ��~[�s���}[,jtK�u<9�*s9C���Erl�1�#�R�W6�#��LD�c���1��%c��)a[9�7��X��xe;�Z�\��.�d�����(�Z�1���&֓�����t�������gy��G����v�^$�Y��2o�i�I:u΋$�o���bL�[�x��{Mr��[ǯnxo���/j���;'����K�c�J�eϵbELc��3�D{3�?�>�W2�v�C����?*��[�2���k��\r��W��o���O��.��kݲ�4���w�Ub��
ק�/�r�����/c}�2&k���4A�8��#$���]����ݓй�ܪ��$%Bs�c.V�F�]�]Koi<r�ϝO)k7���]���iGo^aE"[���)TbL�)�Fx�,h���\d��
a'[��"�����c����M��)�i���T�~t>�3�p�����=�ޘ�G��L��a2/�W �G�wo����={Gn�F�J��)Q́�{��22۫�ࡓ���'0�6.bvT~�1�R�@�%�[�x�����]��3���t�E��ě(�l.�N�)h�r�9%M ���G�)LB��4�-T]��[2�Q�c��/�e�F�Ɗ���-{CYaFJ�"zY��йq����s��.?kޣ���E����'7�ː7�<ߋ��p]��Ø�69�~ـ2����zڪhL��Uh+�QK���#���6qfO�1��(���� ��<�&��к�Z���	�}75h��W���A�и���5';��|5z�k+4�A�6��w;��!�p�_陈���? �N�N�,@5!Q\8�_�`�����&�¢3fP�V��.tILjz�&ʭ��f7����ފ}	>�圫J��U}�xS�R�"N9\TZ"�_`R���1 ucL[��),�c+s���4�RyO��.���ʼh1U�t�xe�� ݧw�E���c���x
�q��Y���&�ϊHߎ�e��_�/ò�(;����z��l�J�XUʰ���N):�'lnr�fgn>;���׶�^C�T\�g�;�1O�X�S�b(} �<�s��3{�v�_�B��g�A��;g�Fٖ�-.��xy�p
8��<�2�q��갭����6�\d��	����j}�+�  ���pd���Ĺ	��B8�'rK�J*�_��5�t.�)Du����D壇8�T��5j���<q+�����k 2��k�~�;5��A����8��<ês[��hu!b�18���wwAt ])�$�.�V �r��)V!�T�R��,�M8ߖ���0hX{�����3}�����)���!����� o���S���骨sj	3B�� �rƎ��^���λa?�a�6ð1��'h�x~�(�$&�]q����&�DZ�S7��T�������8�Bw�ךZ<2Yo�[�H���~��t5v��	v�@������ȮT	��:��e�/�$���FFb˫����[����4PT���n��!���D,�3v�u?��[�&�0^&�d�}o&x�N4������������r^E,�Q�JD�_�\S���Ġ2���f���<$��G�]�ȕƁ����}�ǲ����U�z�#� (mo-�Q�s괣�D��; Xb]�'4��[ÇX�n.�'e�,9�����ĹB1���(ҲC����̛��V��;=�p"Oqș� �A�7Y0NZ	6BƦ6F����L�7���)<pM���K��P�yJw@�7��H)��o�\�6��Z��K��S����㇣�/1R�9�&�.�/twY��_Q�~1�v}C�|W ��$!��4�+���Mc$���'1T(���3�ǽ^�vD�kN�9��������B��c&9�ó���+c�J�}�&��]�@�W�a	����O��w��a�(C��w�w���Sv¹������kh�˘雘��NI#�Jr�h�RV�p|�ԗH9v�A.��g�'m�5I�����^�D~��)C��G&�8��b�s:�,�0��J������`.�)L��E��� ʓ�HB���Ar�ڵ:p��G����^�?��y\|Ж�z�;�؎����aB�}���2��PJ��bژ�a)z��'��o�ۓ��^~�G�8�{d(W��J\�ⷹ��`���%Qw�`P4����2�Z;���(q��J�C��=p�h����@�wQ_�/{q�m������q���f�.2��8=��~9�Ca���nK w�����c�aI�YO(��NL�Y�$��AM��A"��(��CH��kF�&V���	C���Ŷe�"�Obء��`ҍg]�e��ԀQ)4�Sn� ��F�LV2��bϦB������2(`x�1�w�ڬ=v�q�;��oz�mC��/;�	�a��*ki�}��m�>}FDd����}�_�g����U�ʯ���2��Ӱ�5���(�EB$Gk^�sS�Q�E֓�yWÈ�6�obo�7�t3̋\����U�O��L[���ʨ���AfIVL���������C��_c��sM�Z�9K�<FV]���ӒPߓH��p��kJ�*�u���"��G11ñ��`V���갵+<��m��>O궜�6A�'mE�L�\d3����(o��,���SS"��4��X�h{��TǾOx�P�u��>�������&�P���@�����s�q���
9p'�@�T�t,Z���U�B���:�??lܮ�3!V&�>IO�Ċk�o����2��o\y˷�-�� Y��2$+�>�󻄄��v���il��%axt�=Z�^�!�B�b65�>LĎ8���E� P[q��*��O)>��j�opգ_����nQ�&�P!F�$�;+����������ւ�G�l���^t��_k�S�K8�ቸ�[n4�݁�%1�@�)�V�92D���>�m�d�Ƈ��V>� �����ͽri��줧��Y�J�qs�(�z�s:��`[�#ʋ���8�i���=��PK��CY�I���?�.^6\L݁��@�����9���Zl�`��E�P5��-�2�V��Eo��׀#��mh��g�Nd�k4�%�k8��i#�״\1j,I�L7W�d�*�@�.�wZ�08��;�@R�cD��#��Ψe��OJ��X{�(l(i�;��#r�k��(aI��l� �+��l��+�*��'<�S+�2��>U?ƨY���3M}�Mz5��G}���"10)#��cy�C��5��"�3>21�ʧ�����d�ٖ������K��8�)�o�j��
��x*�Su�KENǫb�/.�c wE���=����oHV�jG��uj�5�=���$�,��Oj���/��D�E-v$��]���c�� a��,�ۓ �&��{����P����>�����`+�#�cY�al���<���l�.N#e��}@�Զ����r*g:���ܲV��_"@<���Oӂp����l�悈���X�"{;C�Zb�z����������V��KCM�b�8�� k��Q}���ڤ���K+��1�'o�!�Fs$����6!��nZi�s]�;MM@� "D�"�D��H��tN������pJ��=#m�c��;�XѬOC���(-Y,��AJ��|��=
������7T���3U�39�%��r�?�����W�_���������|2cN�mkZ��`,)C:�?�&7r��(���+˴˸��;���.�_�tU!�L��F�_��X��Dz��D�I�&�|d��I�a'N0&�q��0���R��S� ����s��a�r�W�A�~�� �գ�)v\F�myz�?�*�A(= ^ݝ~V&(��$���8�^��O��*�9���	g��)ӏ�Ggz�ER�A���|�ppi|���@��a�"�<U��J���B1����"��/��pkj�|p�cX�lk��+�3���n�L��n�����^��c��#/@!���xɇ���4��l�ch4Zn��9�M���X9�́��?���������a�t8ðIQ�=��A���_����5Qr�!d�|uL�s�UZ��Ά�o�d�c`fvR���OB��i�`tR�(��;��q��T��_2P$o����6�.���	��M
A�+�_��AڙQZ`�ld�X40�^U�E�ĭ�0mG߬�]�_��	�_�:mN�w�S\�2�m��WI0\�k&�������y�S}<��uPUU��y4c���lHM7;+L]��u� ����f,d}�:�A���B�`b�fRs"2����Ä�1PN⠀�`�������5��/�>&���놚�(���^j�o��>���8<�T�i]���[,��a{%Y w�F�~5Z
��d������-
28���/�j�F���4t����s8|"���]Z�_}������D ����}bXu��p��|j���<�ܒ���h��H�=	�Ǟ�JQ�[^�|f`��Zq��bZD��c\C�Z���W��ajj88�h�}Kp�nM[1��_����j+$g�ԗ�j�&W�rUT$\%�5i�0n>�S��T���u]-G��]�^TLC<a�[�N�	ϝK�I-�����q>���W���Iv���;O}�c�@H1,��&?x">ʮ�]�Ya������݆�a�>7�=�i�9��U�Y�x�8ir	w�d$�s���e�\U$�^������rm��n
9I

��'�y������OK��/%����2#��	�����Ѱ]QV>�����薆@��V���V��{ui.�PR�����q�bl����	��AqJ���V����I`0���y�iެ��e>���M�Z�PAZ�g��L8I��Ȋ�o��b�(�LG��U�~;o|jL�"�@�=�~{;i����m��Ƣ�Eo��H�DrV�o�埜F��Fh	�i�>\`���j'�R�+���l��)�}[�ح S���zDR�0
�}��ME�u��p,�7�(���,�����G�}�,\$3�x��|��� &,�g>gl��t��3�m3-B��0�#|��L�Q��1LF.-��#�%�TT�M�V|`t��rc�T�y�����+6�$��şY/��?�'��Zu)]&Az������x���uI�X�;|�4(6LTL�{��d�c��L5������"¾8�.?v�� 	+\� ����χK��߃�W�����6�[)���:Ak7�	=/^�������s��o!�TZ�X��E���-Q��'�B:��]��_2��٭���g�~�:I7��E�?f�K���yQH
:O���%Pش*� _�����v�����>�.>!��:z3R��}=�gq�ੴs��`�P�W�jY�M�J�ic��%��!��e����]bS�IY���M9�� /��]y��f��F��{�l�YH�ϗ�9��@��@��<uj��餀Y_�>��8�v�S vWj�lo��so��i��\3D���&�!�2�>K#`b
�v��~�%a��w�ݥ�&7>6��� w��RP�ؓa�hZK�U�!�c�ö0{�Quu3z�h0�/����H�Glw��Ϫ*�կ������<X�z)p�riU�M��L؍���(�:�O�m�{#D�	+�� ���^d�]m$��h`1?��T����]f�"��{@n?g'��Ў"��RU?K=���o��d��տ"����C���&I�E_������H��=��߿H�Q��:sYX�O�%*\5�~6�rMq�!<�&��
|�'�i0����^�S������\���}p�&�J���L�
�Cߚ�F:��6A�T��F��rUQpv����bN�C�M��"'�Aw�񽜔g��S��OۓU���@ZѴ�i�F�:CR\���"H_;ʹou��̾<y�����P���O���靿���Q-�'�uLg�G߫+�
���P^�,���Ԯ{�r8CBz'����ֆme_`�Uܔa�B!��'�C>O��7����J:~=�4�U]�>�W��d�����ų�>�|�a��nX�����f�x��A��fs�̮�W���8p���I�������
��pD��*Y���-L>�[-�2R8x��<��j�ۻ/�M#�~�T�O8�`��;����gR�{Ï�n�W�� L�:ʛ3��#��L{?-�٢��(o��Nv kϷ9|F<�Y=n}�ػ�/��i+̰f�Ɠ656��(;�z�o����F(�?F�W:�y~��z�ui_V��Q�&l9�	��/�՜O�jI�)��0��ԍW>DA7�{���)�)L�ړ]����k0���LlRXSwͳ����d�(vi e���Ew}�=��L'�|~��u�[�I��յI$ ��$f0�y���mq㴦b�C��ʠ��L{�^�thKvNLo徇v_3�}19.�]
=+���,]��h�}�:D[ ��&�Om���QО	��rٝD5���k.I��A�958��;V"��ϑ�P�[��������$�We�a��9��_^�>�iZ��΄.����!����W�
r�♡X"����y������(�ə�:�3�!$6Rim��,M�J�R�`�o�r��R��*��c��k����h�S�KZG4�|��e4��9.��/ 3 k�/�� w>���l�#p{�L}�}�Kƣ��0���������(����L�O�R��CV���.�6{�A�Ø���R��Е����1�����>�����y��n*���1
q{�og�>mv�6�Ц(o�s�xcn�`����a��np9�����8(�����FF �*.1�!!����51e5��l�-b?C��l�z�)���=��G�t=4j�1`�2�=�b�#E��C'���F�75=�.�XQ����սB�;o�P.q�y;�Kc,w�5�7���]�)��,1*1QJ�~O��<�'_�� ��e9*�a"�>a����9d��@��d^b?r�8�8��.�`�Q�Y'2�4/uG��o\�+?b�Q�.8D4��R ���"^)�`�?�(��3(Gq����ז�{���,~��d�1�K���8_MCE�8�,��ІN��~B����U����G�Dfy��07T���ޣ��}�o=߫A2�#��j�rc�>�K��i��f�:}�Ǵ�d��T9�M�u#�W��qk�U������2qb��4�0�,2�\.k%Ek-{��B��V�N�R<�����z7�h�V?�\A�65<�C�D��-�ɰ���0`��j�gg�������l�r܆K���Qmx������[�����u/���Q�������&�A�:��r��~i�����x�+�L�%>�t�-�1�z���ܿs`���l����m;
=�~�n��7���]�h�c�K��os��bL���U�>�ښ�F��˞G@� /�4s�
0K�њ��@�0�����~��T%�G���A�+p7��j�������_�--+�k��2U:vΑ3If ��7&\~y? �ԋ�pB����7��KLH�BD���j��{�C���/��Nx�;�ʣ�����W�4;���<:w���̀1�Wu��:X�cz�T�hJ��R� wbz��.�D����F����~�|a��oY c�v��� ��rgp����X���<�q���O[VzN	�"����~">~w���T�����iztGNn�N������/����5�aŹ紘7@�Z�pZh�k��J�Z;4��ݰo��Z��~mS�X�S�
��:���ؠ�w���ߗ��g�\.������V\��5����XH���n�[Se�'��WI��Ծ�X�����!� U|%�����/�������!r��噋��ڈJ5��I�+��V�s�9ؒ�b�O��ڌ�Ӽ��y�LfS���)<{��<�L5������wh��Yυ���;�|jb�wPk�!mh��lV'~ӱ�X&-�i����_�|���ḳ��d��ݟ:I˂�l
��י5>a���S5'�-6H�c8X�x��S}���S:+��}�QB����v@w-��r�k]�GŰ��.���K�[Uh���m�	L3;,P��b���p��8o��DM�
� g,�́�
ܛ.��Y�:�G�����P�l������'��}h<� �rz����=�?�+�<�٭OZ�Pnia�ޕ�8^�:�0'�^UuA�)��H<�WLMN}����*��R��{�П����ޑʛ�(U�'���-(�^a�߯&��x��j>�}]S��У,J ���엕���z�0�d�<b�`� �����4�X�O�_��,��#ߩ�$T��������
˔���Ax�vF[ӕZNA�(5�sz�EB�E���r�K�>�U�>�fǬO����v`ɲ~f�S���uz�	X=�;n��$�_=�+"����=���`�1/�eI���Phb���7�W�3K����y�+_���ѧD�Y�^�S&U��:�����%������փ�͔���I�ԛw�ߣy8e�7&��@Ⱦ�M�DϚ,�;��g*E�P�I�����ļ�2���r~�$��:L�I����S�o�����l"0A;��cI�h�M�l�_���M���8�I��H�Q��|��b�Ҥ��v��	5-��>�3K=��r=aG���Lz�2Xo��)��+�$�M���V�����r��d�w�� �)�\3Uٽ���:���}�V��P��M�d�.^�Ion�P��Ї�b��҇NF�W���~������̗�M~�<�/ٰNZ�K�>I+*Z�#��6�d4A���4X|��s��!������ǔ�hG�k/w@;�68`2Lã�U;�p�A��ܳ@��Z��'T�j�E��ȟ'ן	'vɥW�#/�O�H��r��,fEn�`u�@��%�� ͍�Ǩ�CK%�񉐘G���ETL9�]������X_�����Umh��a�L�_����'��Z���+�h�Q�r눏ܸ�im	2
�U^g�+�B{8*�&�G��V
���!lܥ�x�?�ݮ߅�����|PJ(��L����nv;��t�� έAx:��8�&�е�������9{�n5!輯5���G����#waf��k�Z�%��z�#"	�7g"� �`~؂�+3ʜq6�HSQr�)�u����&B����|�ۿJ˾�eǘ�~��E��ݑ�/��l� ��?%L������.l�X�d7�x�R)�V����$�s��M����́*:�_���"�������2(c��@*@P��Ō�Q�ó��ʢ�n+����1�9o�+ҏ�Ak7�h|28>�r�D�QtYkq��k%�?q7� �,��gpJ�Dգ-=�O�<۩[�w�0/�[Mdb&��������3�œ�}�w���)|j;���C=o�@�B��u�*�=�V�1ÁF=}�2o vAE��L{���:£1iJSBcI��H<��+F��lA��z��F��tq�*�P��5Tq���T�U�����Y�BP$r �ؔ����������
�՜��'b�1P۝l�����)��w����+tB�!�c�s�h8ll�<�>�º���!��	QΠ�1,?��Q+�@�c9>i��n�+� �|�H8�> DcHgy6t1�*p��E[ܺ��	
Qe��>�7&]9ԭ�T�>�ص9,��r���;¬6�U|�����W ����q����m��=�����C���5��l�ŘqDt��)I��N�6싧�������u]V?}�%�I~oten���Xʹ��/$��ѭ�3������rI�DD��'~��=eCڽ�mFs����_���H	V�g�63]���=H(m�Z�K�S��ڦdd��Do[[��Sl�4 0��$�90�_�ʄd{ܗ{u����ţ��8Bg
%�,��Hc�ׯqХ�s��B��q��Nq���!�%Au�r+bɀ�J�"���Vr
�R�|�gW��'q��"�+oR�\�E������R�?9̑>�D?m������mD�D��d"�}�+PeH���.Q#��N�s�aB2Rʌ����Q@��F���:���VG��4���K
y�[�
�^�^������6m@�5��'d���ɡ��;!�}�F *���Y/�`�>�������xߔ�s��\�4�`L�M2�8@WZ��|O�ۖ�`�-
��~�=82��ϐNw�Q:�����[6a��'/Sc�e�	8�`a��v�����c�Θ9 Ry�#;�����~��_����ȃ9J�������ou{D��,�rR[k���5��-�?���&o�m��#9���"���a�`��z	<��WHyi+�c���	���I��.�
!q��+T�ٞ�!i׺;r 
�	�\٣�2O4���tV$U?��Yds$�g=���e"K���_�'�C!�3�����8�j���y�̪�:^�oYSBUђ@͊Qb��\7��h��b3��k���Ee���W^<F���w6��X�W>�ϧ��F��j��o����
�&�?�Hg���Z}���P��Z������K��E�B����e��Y��:�|u2j�Մk ��i�f4NJԔZ`�W��P�����(:%��ܗ�)P�,�r�x^��J����F�w���	�1a$^(7���d��hWk�z`k��6M}��NL���;��vd��)�Y�7�w��]�ɪ�mj�����:��ν%����R�V�7�J��������'�̂�.#�Fa�m`^����i�����xʠ�=��v��(�cr�G�uf���T{%�/�~s��a�d��GY6�Ӂ4�b���,\�$��>��t2<�kJ~�Z#��G���؂�݊&e`���O`ӉnjH�XXJ}�5�)�"�j;�P^���˽Vx�yo7:���x�,zd	����7��l���9;������)�o�R(�2���ꑊ"�y����X�5����"ܱ���ce�jX�Wbq����g>����v*0��|�K9B!����w9���e�w�B�V�ҩ�U-0&Db���w������:�����|x�����ѻH�51y�����Z��ge��aq�hί\.��V��X�#��&�`����S�'@#{��n AgU���I������*�ٳ�q�����ӄ�\x���5�]�\P!��4\}�/�,�o�>-0E&�'��W�lb/��j�3����>`�X���pM~��ÿ��f���nL�()P}�����{B���� ny@�1��Lx{x�30�Tg,�"4%1Oix�o�2�-8=�p���S��zE��XP�^M���)KB�b����GWUԁ���w&��ʩ�{��zó���t��O��d����*�U9!} �wNx���|��)XT#�s�Z�/�$s��e�I}�5�[{ZF��mF�ը	=b�阠o������� 3ȶFa�C.aj�<�����0�iפUEM�gm����؃�0AY���9�v��n��������f�G�#y�U����_�_�*ԣ-Jˢ��vD�Y8-�{��Ϸ�ۼ��f�!J���ۏS�kM�;�N�jCM����}�Րq��蕎0��U�T٤�_�2��9��^Uu��S�� �d&I���� �o)�C�k�l�[+7z�Oz$g,�l��q�PA$�;��<xC9�RIz�!������������]^�0]O�����Z�)ܛ=Ʃ�/75U���b�e�K~Ժ��!;����RV0�����e���;����������G�^�f��TL��il��r�jU�QH�Jlc��Y� �'��Bp3��R��6On���'�n"�h�?%�l 9ɣA@7�m,��7�)W~�$���\�S�@|�z�s���A���n5��Cѡ��.��v�l�X>�DKM�G�Yl9
EQ� ���Kp��.��닚�Zݝ���s�N�@~p�	op21���p�F��1�+ f�^-���<�D����C�b������ƨ���l1 �����Y�?*�j|�_�v-�}�H��~��;�ˉ�a?��TQ��t��Ht�ǚ���V�ɩN��0�3տ�y��r[������yom5���L<\�H��U˥��:����ѣz+�z�� ���'��\��`9A.OO�D�y�\%̞��#~�>I���e����7����6��ek]ƣB]]H��AT1��L-l�-��'�R�fz��CU"�����)%	�����3�s�,y���R�K�F0��O����n+Y�� �Ux����qڒa.�B���-⾵1m�Lѿ�b��gT]F��fW�ʹOJ�U�j�Sm�:Ã��*�m�r��@�t�4�a�L��2	�-ov�w_��G�T�L:�s5,���4�Ng��U��Փg�<��K���@�:8�q+:�x���95��������d��bB�*�G�i7�zr��×���T.u�/c71aˤZ�߱���B'2è&�X#������R��?M턭��[d��05f��h_IJ� B'�l;��d��QLܩN�*H��Mep��U��SEp�����|Q���䍥w4��ƾ�:��!�!��lq.�n�2
����L3N( l����T��ΑiE���:��k�'@���; ��]��JLo$T�2=�=(�%����]�����^y{�9�Zұ�Y�뭟j=��<I�k����¥�_�(�~J��d[�9g��V����!��ft�#@�y����*����UP�}D������.��znoʎ_�>���r�gw�'�4�<OV��P��Qǩg���>R_�Fetei�4�4�8�DV<E]ƽO�9�տ�R�h���1:ןo��$���2�N����	���ߝ��C��XQ�,�z�y�!�52�K��|Jjژ�j�G+q�a��-A�`�K�	�.oZ4ĴVH�;��y���槑��h�XH�e7�.���w�������>�ʸ!A=(�%�IkBU�y�a$_E&p(����j��g�e~F�d�;‱��������NÖ^_z;D���:dT&n����n�-���m�;.P�V�n�X+�3�H&�$(���4`�ٛ���[��m���m�k����$2;��v�R�2���g���.��O����}���<R��nQ}�J��d�w�fZ��s#�|���B�ϑ_��
4��,jS�hجZh��M[�~.�c���H%ؽ�n�v�I�S�H���NFa��%mUy�o(�P`r��Iq�C\��{�-Ӟbhu'=��;F��k�Doǘh��*��ɡ��BxK#�����iI����Bϫ�:v_d��h'����:�F�p!�q/3-	�����^�a�̖.f��m#6�/,�1���D���Ć�����9L+ڹɇ�MɎ�V�	�~_�>�:Ya�_#�s���IW1���9�9vfB �LxN2|Mk��ϊI����� |^޼px���(ޒ����yyn�+'$�j(�^i>���4!����D��;�K�\kҍ�YS���`J�&��_Rs2DB���3m���I�-��̝_�I��7<Fm���[;M��K��U�Z��6�{6#őJ~ynB#	bO��u��e V<fLM`��~���{������It��%Q�[�D+𐾓j�J`������j��S��to��t��*�L#�Y$9�YGAF��P���ރ���-�)�(eY��O�(��Z�S�]���zM�S9�Y[Ş�s�V*`|� ��U��e/��� ����D��m�@��g�r��	�#�LM�8�#����Ԗ ���b ����6��T�rD�#?fpY��f���m�B���o0��cܤ�ms��M����� �c�����du�l��@!����N��99�ϐOJ�ߕ������f�k[�5�q.Uo"wnЮ0J�/P��a�tv���1*�������t	��IA0I�50~ŖW�k
�����ѕ�_2i8'X�T\�����UN5���r�NK���c/m�v� ~�DL�TI����]T����|nt��(��6T�_����&�������9����v9\�G�ӷҴ]���ND���a������ζm��V1�%�و�MC�$d)oʤ��<��}?�3i�P�Ǜ�vIs��5��扚�5�v��j�Z^����\p��d��\8��\���ư,c��`d�w���w��/-�7��@4���M�l�<�����&�\�A���iH�Lr�v��LۆQ�9ԉ*��OMY R���`��nS�xF���P?��0�̷�J�m���.��F3l����d��3�9��^��]0��M��Qꨈ���_e��g�K@�UxzK�g���H��o�bT	(>�}I�F�j�_��P��_�w6�mZ]-��`���$O,��.��XR��)����}W�]iLnMb�N��Y	����#_3�CoTĦ��?�N�$�_�M��zǮ��I���2U9)�^���� ��0v��;��;#ueľ��.�|�{�}Ć~��;������_�"�!O�b���Aטb���o,�X�W|f����G+�'���F�:�2��g[�!�����$�	��ݻrbv}�L⸓�K"�g�K�y'E�ȑ���hn����
��R���U٘�P��e��WU�W;�����6���� �z����ƀ��a��o�?�Õ|���%�t����|(30�q؝�P���A����b����|�||G����r2#������q��L�>[�C"��q���*��M���t�c��E��,�&�vG&�%c]P*�W��܉�g�I�-���)�] |o/���.�X��%jNy\I�=��1
�bB�c괇��	(��,#���Mé���U^[�J�̿N+̪�O��eLm����H�:�E�/����]1�#��^<#6�a�N9��>��B�.�ۅO�����v1�h��K�4.���IU1f\0S�n�M�/+E�
���o���l�P
=J����R�,�A�`���;Eq��J!��\��&%���KA	��A�����k�ܺ��	��4@;˂��~m�{��(\T�\�����/u���;N�P�S�S��X�F�=+��2&k�N����g#��gL[(=�Iu��O�f�t	�_u�\�T��p�|���)B^O��L2��>���F�P���
�6~d�A��h�!>�ϩ[�ٵVOW߉M���St���2MP���@��ej�e#��a��F����er�{'�}�x�8�1��a���q�A"O��6�
ޢ�� )�|�����ė1@q�S�y؋5�� �yf��5	B}#�R��u�u����z(V�Ωs������S\Z�*� b`�s7�����K�_��´���D�n�J����C�{9�y^>�� z�'BR����(R��DJ8�~�9��&ˀO���T��7֜�K��
�'՞Q����ϴ���?���߇�*(���ڗ���t����DI�3}Q�WF�G?���'��¸o���~/⥰IT��L9t������A�~o��ޥ�d< ��{d]�`��z�t��e���!Bb��Z�u�����aڲ�X#��,��DJS_?x��O(�~G?V,Jş$	+xq�R�7�!�V��jÎU�R�]l;�ˉ/��!������jOd��M���p�C77u@��V9���/��v$���yn�,��v>����'d�I=-F��S�а�g��x��@-�l,h!�1���Ʈf_G�'��0����/���8Υ�R�[�l�3�E�#�'�z����Ѯ̱=�<T�Y������'%-"��qwA��^n��ey�6����N����	�:u����V
�B�8�Q�%�"�ըQF���� ���D�Q%JrF���o�&�U�3�>�B*���)���q1X����+��f�<>�+8���_I��j����olU���-/Ǡ5T4��r4�a,���d� n22I�%B���CM9`�6ͩ�;�־K1��Ƥmk�|:5����?��r�٫=[2�t���Ұ.�O
<9��Ab����-�.�rk���݋�&��*1,\C�~Jd��8a��5�m�k-`�"�GV�ߣ���X�>�x�����]jh���Ź��!ȇ��Ѫd-���L��G��e�|�b��bmP7|������:���y�(;�$ֲ�Z���!��ĥ�J�|
�u ����'%�z�ʷwƮ�v�_H�������(�vo�,F��d���Og���E��pZ��z����$y����F��i��v��5P���-��%�J�<u�&l��ݖ�����
䖘X�d��l�-�O)���m�����G��[�͸����Z�����#�0��4ªh������]�3��[2��,�����9�vq�n�cz(gi�;L���1�7��(�Ҧi�f��I�����A"La|����=d���P<ɒJ@�� WP��	` N�3��C#B�B�о���8����!����0���K�Ͽj��x1ʀ`Ȍ�@�������Y{���0>r7y����g����țz��� &��;���mV��үb*�R��	����A��{
A��n��坝��#��R�E�;�T�޸`�*���v��`P�U��pf"i�;r����1���ˇ�*A�sUHu��t�cϵoi^-=6Q(��'�T�
�R�ռ��J	�_���6B���*�Έ���(�A�?$WgGUpK.`:Ģ]<�p8KXT�>����s�+q��\�%��s>q�ύ����'��a���+y�F�����^�P	���JnQX]�Zr�R0~Dz_o:ܲ]����@�{�C�-���`a���=ѣ#h�.;n�j�]�����%�.��9ڧ�a��N<a(d����d��.~��5W�#2���,��{|�B�����N�~[�S�b��6)�N诪� �
$e��r�dK�;ݾ��=�)��[�t�S������m��<���N֞r�7#�U�!�S�3i�¦�g���8�:ej�m�B;qp`d]���y0�����ZjJ�}mڱ��!��@|a�=>��:E� ����~RS����8ibX�
�𿏖}2XL��X-\����`�;~�����Ei�n�O"�؋���B� w̬x/dfAr�$��ǐ�t�w��t�gh�g?;/Av�a��kT����o��ɒo����!k�
�z�F�W��O�"3@�i�^��ϳA���й����\�{"��M�0��Z l� ��v%7}��ͨ4HR���Ѵr��4Bc=GeVp5��@�t1c�yt=d{�|D�lJf�d
�6
_��i���5)���k�o���ѥ{u���E|s8��w�{K��T�	=��Cm�%|���ƥ ��G��!��@N-*(��a������ :w��w���z���G��99�/�>9�{f��M%�&"��ZV�'�4�g\�����7��)+)�[�i]Y]mJ�Z��������l�k]�un/��$�3����gHƶM�"@�`�am�ۃ|jur���G҉0�ݜ���#Џ	xc���T0����rQ�Dr@p���dK��S��gkZރ�bg/W>)��ha�6�yO�eiI:�����(���L��Zm�\~ʴ^�>��᧐�]�η" ��qD��0"O^���d�?|�c�����5� �j���:��C
�����Ac�eW,��/Nyś$�7��A�k�Y֤���	׸��X�֝V���C�Hɢs�_u�A#ϫ4c�j�����a�.�<-���\��,��}2��;\���5_��4�zo]mO >2�ÿUt�O�e���?��G��Q�Ղ�C�k�`��Cm��1�.���XXp�ě�&1�\���
"
;O�r���>��f�D+��1@q�m�u�Q�� β�[�aX1��2â>=�(g��)T~_`�Z�o#&���v��}B����&��
Sǰ4�
��MPF�����cJ�(�$�Y�V&~?���O�Iꃲ�Q���D( ��1�O��$��V1��zzCu���zoc�3:�P-H5�?7JM$���_���*����j��W1#BRU4��Eu�ڼ})!?��E� nu�[u��(Ps@&�J�K�[L�'�V��Ni���lf�K��/���KTY�Ś%��*�3QBjs�C�=y3 O=�����NUy]��N֓_rB�7`{Dr��<0)f��|'������Kֱ�a��>M��|��cM�4�0QYŕ����9?F{P)9�و,�kޢ�Yi�h�6��B�4=5���G�6u�H��
�")��'�G��B�EeN'_,0�>\񾽄�4�?#u���A�� ���;k�g����z�١�J4�>[�#D�0^��J?�A9vC톱�����5����@���N�O�/R��;I���V�~q�S���2�����l9_L�:��s��D�����
����L�׼Y�'{��Α�
�@�b������;�5HW�GD	��s��J�	�g4�IP>�h�i��:(߁�>,8�y�a,�������%/z�|H��0����R���|+��MpXj�
](X���t��#K	������[��-ߎ���D���H��[ ��G�W���&C
�z?�Zay�C,d�C��^��r'��"+�P�	t)]����&����a���w�>n͉�W�_�ƚU�@|.�X	��n���7��)ڃ���W'͇H����-f���5	�2��d��:��߀jQ�$��;��,�Y���l��6�!^���<v���6f��u��/�%�!�;T_�8k�(+!�ING��j�D�˪H�8�� 궝/�Zo|ҷ�G.p��]�����H�E5�B������,�&6IQ����Kv�?`j�[��g�㧚X�hۯ���W̽�xP��E����Q����AN�1��ʰ���M0rG#���muɅ��nA(k>�lO���.b�h��h(�2a2�^�y�v�Y^U��j�8o�X��'O;vo��F?���]+9��(h�c�=$x���)!e��xa��S�U[o �ؗdR$8�}�pJ�ͻ��V�i�+�,�xZ3��,qU�pN'�������tXj��]�B�A+,�P�|2��N*��d�V,ƢD�n\ra_���pkP��ei�"��j�~#�[�T��b_�J9��r����E���2�LBٜ�X1%���@�5 ������"P
��|�v��U���G�汧ӂ���g��:+#z����Þ�>��.�����.w���hJd��i,��q5E����!�!�
�����ՑSN'��вG�n�X��K1��A�{��bP�]e��>�Db����ĵ��]#��kѽ UT~=R̂V#A�_�a�7�%'���j��f�7iI��|���{&O��#�H:���AAk^|����^/Ұ��h�+z���F���V_Tґ��TKAR�T+w�|3'/{����r�.s�������h��ʄր���`�"�����E�RC5c�ς>�x=�C��?�Qs�P���$6��<Ǎ]IZ���a.��N͆��^�L�-m��B���u���+�	��y��c
�Dog'^���<�w�*�~h���Gu����~���z���U8��B ������f^�y�y���L��x�6�$E������Rb�ʬޑ�P�P�e����z47�Mf-�ٵ�9�V��ul�(���9E�QV��� ����b���8-�R��n@��M� 9m�������^�;v6��4=��^�uR��9�R��fA>�{ (��^��$�v�L'��>G���w)��D9����Q����!=p�,o���ghS�*�>�m�����n�V��v���O�P�CAU0Ҁ��Ǧ�����]�i
dhá,�MH�-M�T�vu��f�Q��_ͻJ��]h���J�/�P[̬|v������9���h�m����Զ��6�������jK��2�|���02�C�MDn��ē'��,�����(%���k*���b@Y� �Kʮg/�oj��0���Ԇ%EA@��i/�v�~C�`Cի@�)�*����YkV�X�S	8�/_=j�a��/�F4��/Vw�\i�Pә�qx!�����=��:��}g�p���t �c^��j��Kܤ�^ah~��+��CY�3ֽ���v�y~G�{�a�s,��(�%cR�w�q�T�Be�sl1��"�����q:�iqu	���e���Q����F�u��_������#��l�Û��Iߩ����h �֘h)�xc�]6C0�Q5[�X�IٱR3Cxꀺ��^$ޟQ/���8��`�0���JL������͔�����g?w����X{9���r����.،0j	-q��w.�'EQ�`#S>x������� }�p�~C;a�����_j�f1�D�9�v_+C2]�E k�Җ��c˰q�
�F�uQ��̪as�z}�X*w�L�n`��I��/����F6���GU��n�IC�lсz�0�E��|֧����'�F���#��&�����!� �F	�EN���U���\h��;>�s氎[[=8y�>x�L�7r�N�o������)�����;��͋3�;�3�(P�_� �Y��v���ȯ�Mk��� �=���� ��t*��)O�{���|Z��������k�*9/�j��k_�Fm�8������C�,1� ҙݯ������ƭ4I����=|��6`�5�wH�?�L�C�B11w�A�6[orIo}���~	�ڐ�X�H�r���W�L/����lF��r��z����8f�f<�5��.l��	�V�t�0�l~��r�r!T�=�?=��?5��ܧ�H�m*_�<�f��87B������a1~әL���^可��{�| pb[w�J�����d�	q������4���U�ϛ�Wҽ�Q��_?����c��k���W������I�p�g��00�0i��D2�zga	���8R=�~e�N�O��K;�D�^Lӛ2}����	s���9�>��p�ea*�����OqN��->����~�߹��˗�Nc�,&��;��'�����'���qer<T�f��maVi�߆B�i��|��3���60H���>J�p`̏�?�&��n���m�!�I�|Y����o��<�r�k�y��XM2�rG�����_vs8����D�7I�7.��!�K �S�z����ЅA��,n;�2PP�o����͉Y�Y�R/��A�h�ӶS�s�����m ��L��G
��S*�zp[�m��2ۋq��-*���:ZK*p	��Õ�ڔ�߅uɑ��K�m6�d�処]$�rD��+u�֠ځK�c@���K�{��`ZBrEkB�=�aG�jU�7]�q;z�$���
Y�fϲPs�V�+lcА+f�O �Xe�o��M�,J�;���F{��G�m��d�:o��m��q+~��<��͕��Q-B%�\��u�	|Sr�-Z����6�`����5L�P3� 	��q�:Ms�+<6o� 0��gZ�m�V��2�f��W����4&_5+�֖$�p����i���A�Kz�7�[���F-G.��𶦘��[�~|dH����\%&Cq�F����b����O*��D��j�Qsf�T�HG���Ȣ���J�h�=��6"M�c�:�E:��^�1B?��y���s�ڞ'QP�w�A󗱎��ux�o�P��sXIVh�^�F�4���q��kT�:捩��$�HM�_��W0�Z����C9S��!L�/����h?ec�)�u��'
t�@�����$3p�o������YK��i�¦)@Zj�<}��?6B^��p�Zדmb1*ÃY7>5w��JS��bÄ��hIw7z|M�/�]Lr$��M�y��b/jO�٬D��ut�I��1V�Qgr���7<���p�zF���x��Ga������}��jB�����>���hh!۞|g���kHj�<����z��O�I9,�O/� d�6�R��ü�at+.3������.Q�D�+	U�І���Ɵ��P.~��u&e���?���~��f?��v{ �yܟ����B�G��U�V�V(x?�ıU_a��!�W�ly����ܾ��#̼Z�"�eFhHu$��|���َ�tn*�9��UBڽ��m��i ����@��-(%��LpJ,[��G�0����y�h�#�C^�ظ
J����7@I�úxv@qyKh��R9��~w�떇ޣoC1+��Ɖѷi;* G�'ߓ7LF�]���.���ݡ�ᫍ2�n[��=��uB�=G3��f~+�/*������@�`�c��t��R\9�Y��r��u��H�M����[qz�qٓ��H�{�`q�Rh�E��ѭ��S��cx}( �O~��;������Y�_#��4Z��!�e��D�S��Ѵ�)����׊��_�8}��r��ު�2���0�WT�p��ED2�\����3_�rS���ꯊZ�IX����Ј~�ׯ�{������oS���8�A����f�r� \���V;�fR\���3���j��4��i��p��2��n��-�5��[��d}ׯ��aW��$����)������Z���U�j;Q3��0�>�3��1�;�
B�!��,�̦�"E{�����?��Х��v����TՉ��[�?�&���Ж�j6X�lg�*vl���\�
}S,���j�tߐD\e���p��]��8z���K:PԒ%���2q��
��ͤ�@��{H� L��A����ZK����b�^�^Fs��*��E��Y׆5&�!��m����3b��^ȗ����à��	Lrl����ޡ@:��_�GY5�Vl�X���>���L�@5�CJ>������c(��H��Q��T���}�<Zd�o�	��g�J���.��?L�%��T�bC�\0�o8��@!U������R�+�3Q�dxv�*z?���ϗ�/N�br���T�	˒��/|�;�E��n4�|NEo��� �Y��t /?v�Ԫ�M�״�8I�'�����[
�M/;0e�0�*��k4���t+j$.�}�\���3?�f~�+�2��1VS!�_��o�[ӷ��a# J���NNʫ��f��=�3w	�i��`�ږx��~�'�8�z0_IE@���(���?�O*3��T��!P�����^M*��Õ�pDk�I��J�x�����q�1,Ύ��=�z��FC�z1KOZ��Q��l�Z�q�����/�?
�}K$�"��:��H�B�(�e[n��;=�[�?xZ9!z�IK���z�*�
�b�\�/>�%,37?60i�>J�ik��^cs�@I+�ݦ����pS�=0��	}أ�	����� 0y��%I[xdj�z�O�G"����������aH4�e�ASXt��1��M�ښ�w�$^�I<[H�WA�Ԣ;r1ɋ�.2��_�آ~���7����)��G3�a�����(�|�-�}k~םa*�:г�.2���R�ϳ�^��I7�"b�D�8�������|Z����r���CŎ��ҋ��(ʲ�����M�����y�2��AI�WU2�%�_]j|2�d��u�ʭ��-_��=_��4�|��ôs
�i5�d��Kב����S�8����CQ���q��|u+�O��I	t�ey8�.߇5������cP���,>����0F|WCavߛ?A����Sۮa��E�w�H�h@����}����U��k�
A�4N��e��B����<]��Q�
�y��2�7da���#p�+`����,a�X���J���ߏ�㫇C�����s{	�k�A��k�โ�\����@�[���ڷp�6�R�*�׸1�e+��|k��#'`B{XA�CMQB�8�GW�P��cAhH��$�d/[!�-�����gq1R+��D7MOh���`�o��M����b�D���h��w?:��
@�h#����q�3�Ed��g�|ԕ� �:��j���[��>�*���w�8���z�2�K���q�BaWy��r�)߷U�}p7M%+(���S:�(Y�W(Zs5[�_A$��k�ӄ~�isP�I�pY`ᨼ�_�E �����K�YO֞q�\���X�c������2��o4;X}���9 $����e�]���9���kf!;�B��t,���eIC�B@�u��E�/�-���U�,�@�I�
"'ë�ϛ�A�e����%�ݢ�P����f�3L!���u�޾�3��O M|�;C��]���	?�t|N2�k�oY�p2���#�zb�ϥ�w{��b���{���(}0I�K0�>���+D�`�����+��O�Eλ3��3�����-����%��t�C�#��S�y�ϩ�z���Щ�-N��߸�����U~�)���E�@����㗰^&I�t��xEZ^Y��M\��1Ϊ: ���� �u�z~����E���%���P	�A��܅8��$_�77�AX���F̖C��^Ysmj�ɲ�]����L���R_��p�Lx��/fj�e�]�
��	���ite8��U�NO*�A��ޔ\H#;�&`��OWW�n�,�l��g����}���;���أ�71�gқ�{&3�:(�ػr��ǊX� +vQуD������/��yv�-��^��Z��N�채 ke[P�VT�0)LFAoH#������8���#�2�X>�Ɖ� ׯ��H �$���8�E�#�(Vhc%(1�iV;d A6 &d-6ֹ�~���qd�BAdBO�A�WCg�&U0���v��<Md��h�A���"ś���쒱�N���`�$�S.�[yb&FL��xCL#ՐR��*�'"R�&d75QQ(e�Ma �sC�5f��HTI�:qD�4��X�e��b�D�B��:�Q�����ND�1GRJ��qc�8��R���� 3%x�J�oV�1$���4�#2�Ej�c)T�<J��$J6rF�nV��rZ�#q�5j?�"�x��CC#�(g���X#jA,ǩ�Z�V���� ��z2�Lf��R�]���n��jS�#0DQˉ4� ��a���&"��CvH��{�9��4�T���OA$��3,��2+����5j6�G�sl����x �mP����)����.b~���P�`�q,�"( ?;��A�Ԡ�x��q0bP@DӠ��=�%��I�J'�(\�8��f�#���ZF��BN�P�!��8��)�5<R�`�� .ߍ�Q��.$��!?;,�	>��R���i"X�"rk�T���~��DSI�|�#(������"6c�c���t8��Gх��ZF�,1#`cn�"�uosP�����]Ŗ���)�����bR�DŪ�1Dj�z4�ݭ05*��ct����$���Q	h�'�`Q����Q�����d; e#$)h0�嘠��sIAE5`�2�"�S"R�dQ���3M&�Yŷ:�Q��h"*� i@X���<䘙*��)�9,^��cqIdC�6h�V��	C8�����~]��*}lu`L0l�Y@ L��`�]��Q4��)�_@�5�(^�]B�E\��
���.���H�t�B�
L:$j��t�L�w��#�t&U���c��*�SuD=dQ(Q=;���[��H���M6��d�`A8��=7��W��\�RG�[�2}�ǃ�T��Į#pH��	�|����H�����`����dR�?��d)��sk��T������iA���;��(���B�����
)�0{L2
5`5�>T�Ұ��������Z��Q����)A��)e�	\{�g49��*�����`9���$�i*��@�\*���7ԪP��Atx���u	�!á$�2#(aK)� ,Y�G���b'2����B��Z�`�ސ�(���l����]&yP�p��N���zM22[�z�J���Ȉ$Fp�eGmX Ȉ:C$�k�1�@"����LȄ�!99�4��8�Bi:��#� 3�S)"x�4�VR\�P*��D[O�K@���J$>;O+6
xz��δs)F	Y�F~�f�H&����S�t+Btj|�J���nY�T`� -�!������	hL7���$�8"  )q$/�9�b=���3T|,e��Q��A�ˇZ�J�A���� ]��s�#���S��+.�dFV ��B�bdj"˪R#hr��$-��1������<��1!	�蓮 �ٍ�鰜d���"���TJ�r�F�1�S  ��p!(�FwjͰR���b��l��(!���0rF���amȠ����X���2��i	�t�G�1Qe����#��aq���2�AKjl�FG�<.�o`��9/j�:3�hQ�`9��� -�,W���AD��2�=��H�̮"$L���2`��X�A�I��%��.	qEY�j�jEb>����^	�'��|7�T'(3ǔ0�q<�	��&�U�9�@Pñp��0,��e�)Aƹ!"	��Z�`��n���J� ��"���&IMVc�Po��y:�8�V@e�2��Bf���_��(U��Z<6�y�	��5a�AkwѢ ���x���5(/�� B-�AaC8�+ł&�5(�1�8���q$Ў7s=A�k'q5bא��:�c�xV*�d� P�yHDT�$�t\T�xb{�9l|�"̗ t*B��C� 
�O�UQ�r2^�aY���H x�0 �(�49.�mvHC�z����qbV�C�X]0�PK��"6Se�A�Ta�bPmg�i�G�@u4�2Z�N�O�UV�"���V�գ��.�"��I
�T�QL!��q��<�=�Ӊ&"�"��S���t�'�9�j�<q�,�H���T���1�>�r)�PQ�&;��1���|rl��B8�ʧF���E��N���h�n�8�G\N+K��Ќ<�	AGM�|"6_�5��,�$��.;م�S�d/L�� AXd�i�jT��d�ߘ*� V�s�T&$��:�M����aG2*K�eG���|�(����ܢ%����&��Dv�� �|:[���� I"u����#�!x��d5�C�a��Yv��̰YE6J�i�:�I���/�}��	4rӌ2��U���js�a�`�b�zH%)�$�CAAD|�A�{�J�O�9��CR���R�Ge�I�O�R�R�m`s���Hb��x�v���ϲ�Řtl<Cf�� �#�B-Q	#t5� ٠���bԂ���	��!��Ȧ۝�X�j,��Apt�حQ����&��`������.���\AĹ��\�&�R�U��D��l#(t8H:�cEF�Iw�Ũ��Cra,�!$(C�����"n��Slb��*��a�A�<���2��eDf��"j��Y~� ����,-,��
o�,t�m��#P�8a��;h�� O�P*%nB�;f��kc���| �
�6��ϰ��3N�hV��Q�Enw�M+�&�q.Yn��1��ju<�K����I%:\����S�Q�q
��'�`�\��X�����&x,f��3�G�� n;�n�#�ؤ�AB:�ǒ�r!k�
-
<^-����p\-+�a���8�/��@����z(N�P�
�X���z,����5l�a�^����r �#Dd�]4�-la!x*azT*d@�E��)����D���|�<*&E�4�R"�e!=Ie�D!��)�r|J,��d��C�$'N�1ub�\��ݐHđ ���1��A�\�9h��-L�ʌ0da"] 	��\y�Ow�!�VD��(4H@L�0R�V��DpP-��>�VjU�tF������X��B�8��H�(�g�@W��|��� *�e6�ZT$��$�����\:�,ba<F ���`��/�*����9Y�L�Ԣ�� V$�<T���X��D�M�z�41�@n��}_#�(�+ ��Z���Os�U������ZɊ�����`c���l�G�r5R��wag��H<6�ɕ)����Y�F��됐�f�2�� �˦M\��Ê�,
�⸸,����dCT
=��=�ҢB��t�2�RV������ʨR��i��#v-jH���PfTc��a�T+7��愬T���	��h]"��JWjA�Yb$;�T�J9��-�X*��錑���� *��@I��s����*����yi Cɗ�F���c@�Ǌ�D���wH�XR!_�E�TD��R�c�8��'�)�H6��[g��g��I�`v�̉�r?H�B���5�-���TI}4�03�� T��!D�4��%	�RF��P�[0pz��l`�,�����]Tp�*UX���VrKY&+�F�� �2�%	/���a1��`u Q8!���"ƌ�3�D�Â�XAyLE�a�GN���d��a��Ja��0��ۅ1G�%���h�:�)�����5�]ZCqr�uL��t��E�D6LxcV�c�l����1����kФ4�@���q$�=b6��=�`G�|�7*s <?����T9b�ӝX����iq(�#�D�!�2���C7{UL�#lS��dà&N�L���nL*dJ�N�2�dH�4���E�z�"Ɖ�(Jk�UJNXB�4<I`� j���q�b<[�����@�$`Dj�ت�|F���#����q;oT�,N�������U�(��@���dTU��c��kYB��5D)����Xѐ1�]bC^��L�5^%
R�xSHsJ�֤��v.��Ǜ�� �c�,~�H(�㝆X��$�C��VmF�>z�R�
I�ᄌ1�0�ت�+�X��b�$������PG�R#���5��{	��ofK ���$_!��v��U��D�PrC��&I�&/�gIt=C-������Ǳa���u� ���8x����⩈��	S�JP*d�,f�P�4?U!�Gr�Т��"[f��T�^�ؘ.E���X&QiD����M���2���}��N	������a���1F������q3e3����)l^LH��"l��j�Xd|,�D$+P�*����l;V�	�v���3�R�0��DJ0 e�"D���Ƭ��<w�S;�v�&N��1�\%`�j5��,�j"?���E�����&*dvbJ�^��=�{c�xy~'��,���
���� ��{�d�c�qQ�J�t�C&iT��	�1����R����r6��#�B"S��X��D�	�j���� Y�@��h!G��B�O�'��R�%sXh��C�ݡ��%�Ŗ��:�KD�P9t�����:�T��r)t��D``�awp�"�+�8L�ɍ��@��
x2	)�repT˓qe�XU�&�8'+f�� �7�) �m���[�˭�*�J0$W��rI)�]iX�uQ.�u2�|��L2(< ��cj�I"�ih|��G𾀓l
�Q1U�T	��A�i-NB�ߩ�>�P�d	�^������~��6�6�7&?�[l!#��nA�oH�1�>d2 &����ay�f���DE����I\���36��e��d�]i����أ'�U$��g�������FC����aa�'��h�#Fʠ"�L��(����Ɛ`����J��MQ�70�j?d2:�8�ņ"b�	$�LF�V�T>r@#���V�$5ق8�[h�M�Ç
M.3V�6B��|�Vi��b��S�#%�5�)��QȈ/ ���=,S[���y�>�Xc@m�sl
#��2�>��j�>��g�Kpf��<����(KJ	�:����7J���(+%������0�T�׈eG-:�c�2�QM��	(���ᩣt1B�e���UP�-����H�d4�MΥ�Q%�m�0L�t�Qp�4�/°��p��ɂ04��L��Q��2��I#d j~؊X��)׆@7���tB;̑�a��U�d<O��|�@"5EIr�Ҧ���	��a��S�H��UZ%�)d8�a�?̈�9�O�ӱ�.�]��AQX@�*�T�O��~�ΏFh:QB���\POG�d�Q�0�@"!&����/�U��t#z-$3~%�(�.H�v������i�.X��J�ʰ7���l��3/ȴZ�8�R1BP�	�֘�i3Le�"L�;��� ��A�!Bð?j	�B�0�F�P�.���Ő�� ��uY�>��돁�4@&��&�M̈?�W[J
�&�̞�T(���pPlW)�&<Oj�4r�5��R�(�r'^���FSP-�H�i'A���
Ա�L�T�b ��.0�r�T�'*x�P!���$�"b���`L�P�ODf�b�Dd&�ڭ��V��#PI�?6�9T�R$t�e���z�-f) ��̡��B<UB�"[��x�F˨Ǯ�'``5"�2cTU(�:������Z��c�
�0F "�H��7�H$B�B62�J2ؐ�E�?�y�(]§�d���GM���8��.�J`����h�H��:�������}&�K���.4c8A6�C�ȵ\С�۽R����%J��\T������G/�0�T�W��0�"Riq� �tR7`SD�XU���.�Q�t��A�ɂ^�N�"HpT+�Lh��Q,�X�$��˖B<sX`s@BK ��+c�t67DS���
಩2��\!����R����9
��^J�xP�O��P��u3@;�7i����x|"� V���T�!W�$�R�Aǣ7�m~��Qa�(bq��Ǖ��x��.#+��+�L��1��9�t��$�{� 	�y^�Ea�eX1!N�����J3[dggb���d3ix�(�"�a�6�i� T����1!�F�L�_�3�Ш�C����PtZ��#����8b�H�#�V�-A'jsP�n���n�������q��{@{��0�VrJ5C2�c��cX� ��]F����R�8���zH������F���&��,FOXR9�ԍ3�A��I�$����H+��s�VX0��8�"���*X�qrO�0�~%-(*�#"�c�!8��qa�C ��T�/�t"�h�Z�YB���2&	�5	Q ����,b��x��au�bt�c�Q,��$�̢��[m	0�r9��>��RD���93	/ ����8#y�BH*�;Q��!�s]!�DJ�
~�I��a�!@D���98ơ�����n�֤	0A%D�9$�F%[�B�(V.)V;D��p뙠�Ă���Fp���6��d����`���
�7�édf�D�I�Z=S�H0�(��� `URCH%�y]� A���"#M�@40;1����6N��Nl?���րqb�_/�
�n\��qq-b��_O�Xq�-[�~�F�سu�֭[�j�>!�Mێ�;v�оC�N��w�Թ[����ڭG���Ď]z'��Խgb��'i;�U�v�[��٩C�����WA\����Z��o18�e���Z����g��3���Ѣel�mڶk�!���]�Z���o�*���c�Ό�ת[����6=�Ƅ�PO���[ۦ0_HTܩB4��k߫wR��C�1r�L����Xl���*�F������p��@0�D�9s��_���E+V�Z�f���m߱s��={�9z�������.^�\x����wK������W��߼}W����_k�}��QW��w\-��[����3�n��Z�j�*�w\-Z���[�փ�m�3�	F��`��=�˷��.���J4�w��Bz5��wh�������?���	����,�c|����w�K�{���y3�zv��S�)?�x�ŭ��q�����~�B9���S6nް68F'h��XS
ߖ�>�({��`}�܊D��c��G��8Co�4�P����ό�{,����#\�O[v��������:�JR��w���Z�S�hм�>��97�n���k��N������˰f�̱~�����_b)~�x�̐�Θޯ"s[+V^��?�+>�������m^q�Q��XZ��]��_'��ò�Ey���9�����o��X�g���g���/�:%H�^8�l����S�Ÿ�Ou��ﭠ�W����epg���DNY[s�
��1���U�o�W��ǧ�bk*���i����x끉������w�J�V	S��:����u�\8��)�HA����Aт�+�Ϯ]��Wg�j��Lk�5l�帗���ћS��0�^T�����7>JG&N���r?�|�	M>6�_q�6����ϭh�_�H8vo��W�n��Ck�/F_�;��p��Ã3F,=xܭ
5�nI�ԁ�s�&P���'�M��-�;�jے)ݖkG���|�mc�Մ�6۽���	��mOB��-�5�����y^҇)>ã�ݮj�i���-�]����?m�3���ly����ߙ=�I�k��y ���_q�~�������_o��9_�5t5��S�i���I3)X@(�s^l����⪥��5Pz��/{�n��)���y�O�'�����b�l��������r��.$�jCpq۾T��I���}���?�yx7�ƕ	��8_Wͼ�
����,x��bÙ�d-+6 �)�l%+�e6,�4�����#��qo�ۜ�}��_0�F]rq��m��ԖK��7������7CN_�����h5��^�f�z>�?��?C��{Fn~}	a	/�-�L���qf����F\���W�%4�o��}��[��Za��ۅ����=^��DB�=ܔ��v	i�����p��A9�ɫ���E��������WT\3]�)ۥ�6��ab����rc�f�^������=PެQ��mYug�����r���9�n�&t|X�yok򇁃�y}���������q���Cw_�5,�����ݙp^��8��+�����rG�������K*�#j�3��?�,=��vB�$���o��㚵?&��\	��?��S{��5�����8K{�ڥ^���X�(?V��O�����W[�\� �A��(w����|�{��NN��Tܶ�@nے��.g��);uz[4z�Ĺ�_w����/o�?S�ʞԿ���;��_޴}����G�<����4643��'��E��\x���ek�'�y��'˨����t7��&�OyJ�P���o���
�l�U]jб�s�}�dכ�����,��أ���������p(�<>�˪>��Wƽ)�]�h�Qz��_�����-9��~�����t�)���zrꖚ�s�~�o/O�&ת��_1�����46�{�J�p�Z��!k��z�G�Mh�Tun�y[-YGM�7k�M]\wdeh�7��} ��O�y��v�
h���gs��k�V�P�iӯ��M'�WC���	����=�PR�F�����X;J�����FrX8�ϔ�n�蝏�9eG�=�=�]0/o~S�!ʵ�G�F�t�Jx��W\i#��늋I�u�?�ļ��O<��Gg��\�����ո��M���x��s���0b�1Kz�û��fe���]{
V<�n���V��_q}_7S��|����W}���2+n?�yt�p�!��k}
hi����c{�s|U��u���:��%G�4b��}�/�[�<�O�p�3�$��?krok�����T�6����[����Z��:}r����(�ښ��~��l��˞`�'_���﹮�7�!��c��̃�����v��e���S.]��v�L�->��q:�eڱ���F�7�3Sl�6�ӧH�>�ij��1e��~0�o��+e���Ho���c�"��������4��7hx�[H������%>�L�zP6��9a��'���칋&�e�~��>�)!�'9<1w��Y������O*�/ԕ�$�n�x����$�?6�6~_��mƄE�o���%�MK�8�~�@K�P��q��ɍcfs�����&���E�<�"Z�Z'X���ݽtf�&+y���{�������}�-S~��Xj=D�i�E��aO�<ccC �_ւ�>���jc�o��c,E�b*���e�������j꬏�Ż�.^6���������)�����k��ɩ��/���k:\�2�T�4j��Vas�>=�����R��̬�����J��a9n:���mJ��g�����+�/N��X�}[>�k���3���?�����s������X��K~���sb�?��s]p�q��0�M��k?����ǯ�e��+�@��?���e��J_׫�U�-�M�f.2Gg,=�I�z�c���U|I���^;�,r(^q�2�}Z�ڴ�Y�@�:ir������k�jӈ�ݯ%��/&w�����|��帹�����~���X�@I�}��Ν�5=�S����ϭs��m9d2edvv���	�U]j�#�C��lt�~�䷷�����Ζܬ�ryC�#ԭ�|y̛Q�Ɯ��ݘv�A�E�;o��������Y�O�9��,��cϯ�W�ϰ	��I�?wN��n�����h�M�N�2�'\�6���_�<�F�����=If�ْ_`���Q�mo`�������9��xN�,X�%nTڮQ��2ޕ5��I�!#�T���r��*�ˉ�����z����x�TkY݊�;�X0�W�ΗOJ�=a/�{۸����(nO��ސVj���s&��zՉ��틖\0OJ/�e���\|1��ig�a�z�H9�o+KˬZYV�ië^\Dܹ���nx\>���/͡,و���?aϻ�^��?�,�i��7�V eH��5���C�u�7���O�W�.�<1k���'�.]Զ��c��zĤ��)IE6�ػ��OHi`�m�<����)��^_S��my��v����#Ȝ�L���W\�`n�%#T�|N㯸qM#�*�7ܬ����W���Ԓ9N��na^އ\��)s��0{Ӣ��_�������	�u�|�Q��K��u�5����;�\	�[ZG�NNNdtkN�-mt����)�-|�~[���䀿�ԩ�K��w�Ve-<м��o���D��C�b"����Oc��o�	mIk
~;�)����璟1���U$�S�!=���=I�3���_�]C|\��ϙ�u�������5?x����ȸ�)�&W_K�~:�ÜST�L<g�Zq6����%����,��~ŝY��}�x��	����Y]��Y��mkR���#9F��pxӞ3��6�ϻr�^τ����Og]<s�s9:B������֔��O��Pob�����+w��,���G戁�9E�v�ۉ���2��������"�
�QZR��4kl=K�5�:�\��b�ld|�toe�-��?�%��L��#vE��o��V��Lg��+�(�_�0l�L�6c%8��=�j�Z��j$���w�Ou�U�-�t|rF�H$}���������}ܹ�}�X_��!��}z�?iT��&��xW�D�������g��xr����e�z�/IF���ٔ�[��%�oY�ѽo���|��%��5<����ݢ�i���H�D�u�W-&g�����M�?�*�l���٥!�\�	Q�f�C�T���[nͻ�t�JC+��</}t��?���Y�~e�u���t�ȶ������W���n�����oV�����4��H�V�q�o*8Ax��\�#!��x80�s�z���8#�C��B^l���h�|��{O�~��z�����
��:�Y_���BI�j{����?&z�M��^�?;û��c��q�K-3mEy�\�g�8�+�Y3(��4Ry{Ifp���s��&M��6`�M��)��N��奆6������ˊ�i��LέZ����8���d���[����؎�~�Cf���"��ٵ�����;�ME{�{������\���g��UO�>D��bN�)]���5%~΢��+��.�.�f�|�?Vi�l��3T������r���n��c�1����������V�ȟ��T�苢�N���Ս��?)���<s8mk�kf���V?�_��v�]��iGv�|����}{�c�o�A�_w�c���wb�p��k�!�COG<ɽL��|B��*򍹵��Q�]߾+�}�u��M�ђ����!|l&T_;�����"�(��{<��}pn-sB�y����M��/~
��/��?�^�\��Y��1�Iȿgx�\�xg�AE럟{�4���9���o1省W�oz���ܐ�'��n�l�`ޗ<�[n�k��~DϏ~9����V�,��K�o�T��c�rى�ɥ'�������mR���a���|y��]=rHŰ�g�w�-HJ<�O_S�;��ؔ�`��U=����rp���H�*p�w<����aI�1�	�m��<���1}��db�K�3�E�j�ߐ������kn�Fd��,1Fww"tn1m���˞�>�M��+w2�&�>f��i���G�K�*u��4��r�!TT1)yÖaM��I3�����L-�v��^�RV�A���u#_w�G��myfu��(�E��6V~�����:wu�j9���e-
�KZ�������N��)��(w���_mM+����������`[��WKV��x#%��C��vv�J.�[�4K�=.R������/)ضR>��G�N'Mٛ��پO)5W�L��i7��cu��7�h���%u^��>JO��<��Ň��V*���r��%�������Z��,�_oH��>]���ӻ�׶^��c!=y���Z��iG\��3�q��ip�N�I�����l��˦��X����ϐ��3�ʟ9�"_.�%^F��UN���e;�:^u}Ú�;)93�f6X#�/)ծs��v� 1g�dfN���kU_��y�ȝ;�|���M���SP{�\�zH�׽��P��$EŠ��|/�i�|ݵ�iӅ�8�COzv��t��QOi�L�;t#yn���U�n��񗂻�l���Pj���i���*�t�~��")n��==Pp��[���zZ������ߺ�Ih�Oq��ݬ�w���:���2W��h&�Z�4���]�.���8�~T|p�ܚ���.��s�/���r��}:��mc�O)[�6�ō��z2gdҮm���*ȴEh^����π*[F�+W�/����W�Ϻ}ǽa��7����臊�nӷ,Z�'������`+�8R�?�(���P���*�^a��nۿ�P����<��pL�˃T>ۊ�ѱu���=��33\w!e���l�G��Y%�ג㦗?Ux�8��M3�o[�_������.�>9_�3{έ����+�+W�WJ��y՞���]	�Wv��v(&��n��nhhI���r����H��;���ؘg/�q}�gV��2P�c���/�}C���?����	�=�k\8���<��x�Zs�Yސ'G�ק�]��O{Lj��]�$L��%R��>emB��_r+sVu���k;7v��U��[р�u�c���8	��M��Q;���>'*J���W����E���X�=�i�gά��Y���y��l��#�z��LGe�)pt�c֩[�e��8�5�s�����1%�ء�dO��	�KVD�<�Ǹ�`�_*<9�˕�Ggߘ7�j墸��s�̇�٣N]�8m�A����u��~�KmBT��z��J;���TDu�߳��*4)˼����0�W��/90��|p�΄�;��]�N*ߤ]^w�\���ߥbڡ�5���:Կ�\4>�g�dn/���L�Q2cffJՉ-�7�楞^?{����Më3�p����w槭#���U���EЩ^-�f�r�Q/5}q�9q��y��̾�����w��V�|pp�*oFE��i9+:C��.�B�?U�Y��w_�g�5��7��}W��5*��I�7�������u=.|۵p�[8��z ���-е�:�X^�7zT4d��~�Y���޼e]>oJ�����z�+��6j"eF��u�S3�$��:;��%��νi:���H������\��ic�߿yJ����t?ꓩ�>+�x�ye�c����+�Ӟ���:��I�:.�߽�����ƫ<��8��%������Αz���'*R����67/�N�*�P�������������z�u$g%NZ;n衲�Y3E�������';G���M���[����a���ۆ�i�e�У���y�䣽��+�1���l���7��\2��/S�>�y��i��������?��znJ��C	U�F
ov�f^�ػa��ڳg�v�3Q���|_ꂛ�wD�˹����^]6���;2f=�t<���Z��R��{�vo�f<L<�.~V�`��́u�K���+K�hl�T�$3 d\�D@�"�l�f�S�Fkz��Q����v�d��������ʈ'k�%��q���c�_q9k���ߴiԕ��q��6�����s�W�g���5cV�}@J�s������M�׌��y��F39�&4fm�R?ك���I���snX�FJn�m��\}��+.iX����3�!��c뒴��=)?K�b�o�-Dǳ���gg�����;�����-��}���3K��w��t�/Η��КOO�uWD���%/���#���u�����>h�5����7΋�����%�k�= L��n0��66�\��qt^ZU�ꥎY�$}�S��nw��t��G�-S��_�0���tn^j��#�g�?�a�:G[>�vO|���I�F��|\�j��ƿ��m���m��`.>.�w�W��9���ū��S[�pn��j����g-E��{�����-I4{�W߄{�n�+j�mi$3�*�ŉ���ݣ�<{Q����C���k�=ڂy�^��[���K�<z���1�v�91c)��Dy�ח�~���{5^p���q�i\$'=�{[���;�Ѓ1�ٛ�c�;fNG�4�}�o7!M�_}�����G��uI�����p'[�+�gu��=5�i��/�	�-�	��G�ms���ץ���,H8T����
^�O�tfK�NN�Y�℄����.%t�?�K񸎥�ꈪ0O�7��A/��r�gު�pqe������|ryڱ���w��όy�����K;ܝ��)L�8s�����IiWU������Ӊ�3���Q�����U��y}
t۔g�9	���:�x��uV��u���$_�[h�:d|*�����[����&�����Րk�ʂ	���F�
V��60Qv��}�ǼO��������qK�9�{_��λ�-��d�V�kv7����p��E�d1Sse����$H���"7�m�1ze�����]��^L<Wݪ��K&������3Ύ�Y�}�?����wE>����Su���u+k�>֞޹���Dq���C���c���3sr+:=�{��M݁SyK��O�vu_��W��a���qs�ZL���$i��ʹ���'DK�����w�^}u�٥���\������ǭ4w�é]j~ŵѴ#ͱ9~j]�t�k^�Aʒ9y��Ηe�V�Z�p�}9l(z3z�ӊC��j0�V��3�s6?j�׀6����e}+*��#�u�?�fm��s�K��kN\Zu��'0�3�K�q���o��ߎ�Tn�};h�eޑ;3;MM��ޞ�9뺬�=0)�Ι�h>�Zs������"������sǦ��ސ�@�����,�:��hJmܡ:M΂�v8R2�.�XR|�>K�	JO�Ӿ��}[��/��O����(�v�V9��u���£Uߎ��v`�$���B+?�J˫������H[����a�s/7���w�r��hғ�6�g���T��5���.�<j�C�?g�,h<op�Z-�������HH'^	�e0ލ�<qG�&|U�Ip�ER�}P��]��=�|����a"گ�ۧ���i�|W����%�h������y�=Kޝ�����7����K�����bk��� �����N� �CG$Σ���:�\w<�`ό?�v~���:ڥ�ǻ)��K�P%�x��P�Їs��}x�knuy����;��\F)zG)L�V.j�X�3Rۜp����ѧ�ԅS:6X5~k���[�u_�_�S��Ho/T>X]�Y^B���f��õmF�Aq�l�}�M�%|��7��K1��
Gm�z�����Uÿ�]�^ ��Z6��?�W��&�9Q�b�X�tGb�ӹ-�[](+�*�/�Nn�t�(����{l]������e�9�{�N�BWl	����A��%�<��Za�E�o�s�>�l���&��aSyN����ǐ��%��1�C���t:��M�����N�:�]^v�����v�A���I��B���C��į֐K%��ǭ-cP*�F�ۚr���/��Oo�i��O�#h���hQ��� }'����~��S��ѧ��[�^���n`�U��{��3U�Μ�(|m��?j&?(s�vo�����#۹��M��p����]�Ar`�x��������k�ێ�4��MX���ݑ�s?���;+���<5ʂ�C��,���{�����}�i�zh��=@¿ݦ��Us%�v�.댓��kwO�ɥ������5��4��,�Y�eT�� 0��+�s;��	�>�����G#)T#h��� ׼�}����9� ֦Ćo
�@L�\��� L.?i˴�[�c�<m��V}ԡ#;W�{u��:ӛy2C����1��McF�L=�@xn�{� �'�^(M�&�P6~����J��.ܬ�ģk���<W�����G�Nq��ӟ���r�Q#1��=���c�\��X*�Jz6���w��2�z�v:�� .(U�{Ь�yF3�� *C��9>��\dF�#<`���cd����=�+2�3�6^(&��G��/�Z:,c���9 ��k�uI��J�|�ͪy�T��1C�:+\+$cm���ӭ~�~��$���v����'����.��6�@��_�:u�u��3���?Џ�W-E��m7�a� A�d~��ă���x��\���8���C2�9�{�H	Y�/i��I����y>V� xmɓ��?6�D���<1�4��/��+Q��>�2��L�_���<m�p*n�R�:g��,C�:��؁���Z�
٫M&�[��M�����!־3j����A�������
���_���i-�n�0J8��p{W؞�3�<c�MBy2��EP��O$��|[�ZxX�'��˴b7������F�$�rɻ�=���3��1�G�(I%���d�=�<\*����/��Ɔ���_i��0(@�f��E>H��0z��������l\a!ܻ��w&�1�
�����x���g��׊(\~'cU�M�@*��t�Z��eV^�� ~)˚nҪ3�A�F��S��� ?9�o�?J�X�6G���=�X���`t�݅>��ۧ�ՋX����<���C�\�!��z� ���֭C��F!��ߜ���eFo�A\t#5����O�?[_I�k3fE��$r���R��VZN����Px�N[K��n�L4LFA�z�+�G9R;
�'Ğ;��Lo�4���#F�"���A���}M�㖕�K�X.Q�yP���gft�x�$�� Ү�ڽ0T�`�t�W%Ǔ��^M�n�MϨ�  �Z�1 ��[�V��Rj̋�0:q�Q,$�PL�OOZ�H�m�29�EՔc�@��HZ����4ɮ>^Ox��(w'?)8�}sU�H�y� \�4t4r��5��Qx{O�4���>E��M,ڵ�\�K��8�=jψ��|A�=���\�*(Ԭy$�8����S�R�E�F�I���:ԇ;A\��g9l��}iY�����Б���|���$P�~bF)���w*;f��6 ܆��ސ�*��g�C�z~� ���С|�������À[��S� �w 9�u�� �lԂc�	8#9�9�e�I�y��T�x=?�i����N9�:����22{f��q�{P>UǦ1K�=A4q֘ݕ�$��T�!f�o�*5`W�H�^8��@	�;��	�ڽ����<Eh$`rˏā^$��px�\�#�"���;è� �=J�l+>d���Y��>��Ӧ�L���?β�u;yt�N�*�>��+��'�K]P[V�܌�c��-�ON:�z�.>���r���(R��]I�Y�zԱ��G��YG<�5.�}?:���#5 Jb*��W����а�I�''#��kK�@�MI�E�����qR|�
nI�P�Ű	���,q֘�L�;
�>T�<z��W�<v��kS����HQҥ��T����$��k��mtUd*r٬|d��Ԯ��8�(vr�q���W�V�p�@��pk�qE����<;F�dw�q^��!�|y���������Ojiwrb�0Ϯ}�.�_&0��� �y�+��/p�}lF�����K��S�������Q�ֺY�j&���*� 61�t��H7R=9#�Z0g��R��<U�w�Zg��N�Ҹ��+��&�yO�N8 d��:�"����f�p������'��+�x�mV
T7#w^�����g,�f��dɟ��������vyet�1�^)�Ze.Iy��TK`*�O>��� �-r����s�SO�'�9��	�B���"��㹁�@��/��ϑ�¶d���S�
x����;���ۃE�}��H�d��x�G��e���w����x�����v���O�y�~�c_�)wg
Z���&��Q��k�ɸ����vڕ�p+�)� >�7�5١��f�����I�n�^-��������@��]IxX�O�<����2Ok2��d_�ct�sZ��rX�1��9;Y���8���Vڞ����o@6�>���F�9O?z��A�s�$p�ܱ�ZRӴo�e�_��� v�]��Y�0�m'q��?J��>���XL��0#?�>] �ʳ"��B���t��7]��z��]Ŀ	���?�% ��%��?֓�.�qi*�2IS�z������G�5��t{�mWƹeRGݮ���[>[9��%qR«�!Ħ�D*Ai?ʔ�q>���dE���џ�}��L6�l��Q�׊���wү4�6H��tp�n �p}��ܶ�n��Ms���-���F�=�B�G\�u� ��Z1g�G9?ʩ�\F;W'��_z�����H�g�<����ސ0�ؤ�Q^Y�7��x�kԼ_��9���y]�05 �;\%m�+�O�Z��nCy���_Zx��q�8�A����)Y{�g��E�at<������S�~%�Ė-��ic�2�����TP��	���/��ĚZ���Ó�+���� a�~�c����]��I&�����ޔ��?��]�k��fl��������*�Y��ڄ���L� �8 ����=x�G��
`j6px<�w���&��{��ā���׺)>_��:|Y�Ϧ��fp={�Qz���V2I{+�ڲH�n`p2������d��������peQ�ʽU�'�2����+K��u>Q��HX�Q�*4gg}k����v��r�� \���j�~��t����4\���.�q��ԍʂɕ ����j�z��"������Y��~Ķ�6��у�酏�VV�E*̮��<�t�L������_k��.����]���*��0�q���2�z��	�F���םõ4ϐe��1���?¾��]Y��� ���&��ߨ�\t~��vL���,��ꋀi�� < �_W��]&
>�e}0*�� �F��y.��8��N�G�)#�*����25wa��E^ϒ+�W��5W�Zm����j���^��j�ʹ�r1J�=O����O����i��O$�l��1� c�V?�C0^2j�߲N�n�v���:~X�v[���p�2r�з�1�~���,��.$����W���y� f۱d��;�я��\ȾTq�U���s��!c�^�I<3'�}��� _�+�o�� u��V����Q��E+�z����̺��r� � �H���S�F���#���~���+:�-x��i�ס��Q�*el��#^3���|�Ѩ�>�����\=}��V��>������?Z�fϟ~47�[�qPt����'�W��n�� ��x����_�NY�a���0?����?Ds�9�SZ��AU�2�ὅMx�.
�#<b�Zб��c�F#y$U c=sR��<�U�z�T����W:���m�+��@��c�
�đ��-ۮ1SM�<־Ic��R;�P���s��"Eo����kH��>��Ŕ.wp:�$�͆��j���a>\u��
��[���V��� $�@���]�z�+�����¾*���En�J��9���NӽEq�(�F3��Q(�:i�8�ŗ�p�!vR1�{U��ʲ"�wڽ��3j.���'{��$
�[Ʊ&nZꊵ����i{�7(�>���	o#M3��gڻu�n4�A�ݼ��iL7�d|�`�c'��¨ț�ç5jZI���˷��:ӭ2��c��^��C�_G#q���}("��ʘ�Xt���*i����q����ڭ���D8�3`v�Zv�k��H��"��^�wKP��j�$aA��21Zri�e�7�*8��MԴW���A����9�Ul�A�ˏ��cl�+5%$�2Ŝ/i#:��מ�����Hۗ���m�����;{l��`1ޫ�p�\o�Г�E1��mR�P���ޙh��as����s���u������k�kp�@�c��a�1-�zz~�����nP��e�O�Um�Ǵ1�U�y��d\7�J@c�6��#F8`���G5�<�2x�P=W��Ǳ�ɬVybvp��+�~&���w�3&�Y����k9	na�����Y��I!N���� �V�+����^�6Fk:y~Ϭ�B�!%*6�_��fQsk+d.W��́��N?�*]*Ǹy��󚮫��?J �Cn a@�j��yy$�'�z����3���T���{��(B�"ќ��nx3ŉ��{��� ��s�s����^L�p0	���ԼM&�z%�H�+�G�	�U�#�18up��N?,W��G��n~�W���ƍ+�^�m�%�38���x�8���*�'M5���[��Vb�UF:�l:Ŵ�mYT���K��-@�W1�FS���5-k�K�NB�2 A?�y��Gdb�u��5F���������y��� �0�A���&�-߷��J�*�zV�R
���hL�5$��}(�v "B#�)��t��\t��8 t�B�s����/^j�q�\c��s֐��]_�ِ�8Q�Vg�v��g5�0]GW��EoZ�m�Y�0E�w:ִ{M�1��8�^���7�+JYP��M�o�%��Ni���	wj#-lL����y�[���4x�M�/�Y5��!�9���|��7����j���Fc��/
	�aT~-x����N����~�u#&��]�w�ֹ�UVPv���zЦ��qJN�����:��-H�1��m�!L�����V�ƿ'L����ytΦ�*�1��q��� �U����ԭ�r㷮E1F۲X���&P�k�jlh�_����u�qƧ�>���wy1=���U���w����\�����6����;K)����d{p#J�:m�� RI;�_4*,��sX0�E�l���Z6S���O��d�H���:��??�Ғ0\ NGn�犎9��1+�Nq� }>�:�!�B�g���U�%An􉻁��ӥh�Ȑ��鑷��Pl���UZ`c�9 �V������P����������OC���[�'��_2w�V^@<��֓�_�o~�D67�"$r�ds�}¸?�� �D��yj�+%��e�8 ���_���[NԴ��ň��p^�M��~�+*�S������)��%��t�緕dW�^���|҅ �k���?\����L^v=9b>�_sZ0Y<�g��tv:d��F�' ����v�;�.W��Y�-��<�[����f�۰�J�����XXG�X���S(����T"���hlt�J�W��[�6H���V/N*n�mĻf*z����3x�'�d���'�A�z���	W�><��P�e�g%c`��ld�����R~�{h?v��]��Ԋ|�6�t�M7�f�E.>P=���w<�v�7v3��R#8�֗��X I� �� ��9�66��t�/�v�c��qNfܸ^��I��0��!{����[v�N���wpN�9!˩����5Vȁ��*�W~0��k[��9_."G��]��Z����e)$ʳ8��$�)�K�c?J��<�\����HU�m�v>���q��9�R����WQ�x>8@(p= 5�]i��HZD`��5\�V���v@��ԋ'��c�3U#�h8����������� ��DR(�vy� &�ѵ;�����Ѿ��z����d7���꣓ӑR�Ɲ���#�Ujb�m.n$�P���N���;ko�P� i�F�����_����̒�����^������b��E�OlI�\�����6�gپ%���Ͷ��z���>��5�I��0��"�-o�4x�QX�bX�oν���EM�X�^=�3ϵr�-+�h�Rz�'�����T�h�T\n���Ad.��,HV=;���/�$�VPz�isC��1n#p�Yf�q������ȏ9c��^ks�TX[�S660�`���9#��t]�+���o2m �׊�տk�8M�]��@�D�[�O�s��ʎ�Kt
�� �W,�	I3�&�Ċ�|Up.�c�>#'i5���]x�B�P� C'���>������fG�L��.�e�_xSC�K� �7�woZ���6�w����� �\���W�v�,WN�#� c��+�4=b��voq<�Ĝ�ǟJ�f��A�&�l'�ܡ���� o^� �O������Z�Y���_�N@��� 쎦?ޯ@̿��ק�V�rMݟE[��^���Y��GA�iÌߊِ\�ʃ�����n*�<�ɫ��&q�*
���Wm���s�[Ҩ�ʑW���2Y��;O���>��3MCe���%\�z��Vr$�ڼZ��=R�DNZ\�����+��ë0�B�E9���)� ��ʦ�"?����a��-���߷��պ� -��m�ȗ��6�3j��������H�x���r]0	��.����?�f<�����Q��)�&9���xr9>kv���.�O��~��^����ݍ�I����-̻O�~U;m#��o?�\����~8Ă�$Rp?�Mx6��kV�<I:4�-���A�����j^��u_$L���Vs�?L(櫝�[n@��8�巍��P����Ato����"���9,�s�T2\���@M.f#&O��� .�{m�_���EA?( g��y$'�ǐ{�2�|���b�0�J��_C�ykhc-�v�Uq�1���&~ۀ&�7�����xJ8��w������� }ʱ>|FԵ	-�k�� X�z�|ͫ���۽J�7�m;g?�X�^����q���U��<�Ì���\������Nk&Ƒ�����s��8^8�Tmc��"�A��#��?5�,9�&�� $�F���dhƐZ�'��X�3��¾��^�
���N+��y�~��_�y>���d��ӎ��_k��N:���_��k>��ڴ��3V�-G��ϸ�
�.VC�Z��0�3���)@�^U|���Z�O�2q��,�?�0��d��<`�\c��#�������֙�VL�{��7��Ԗ�M|c�F7�`����8� ?�i��<��*}����7���2���ĆC���V��ǉ��f�\�3�#���(�}�c��}���@��x��{W_	,W-����cp ��ֺ�vە违b�6OB�-�U���W��$�<�J�~l�O�I!���RFspH鞔�w9Z��ҩ��ly#�y_��E�Ք��׫�<u�x׏�Y|H������EIr��\m��̠�#)*��y'뎘�y5m"2��?:�@�/��;Q9!5ce�����t5]o�Ê���rj�ڇ<�=kM�4M�H���C����Ĭ퍠d��VV�:��J��It���N�M�:���ŉ�%i�����[1 ����nk8�UVG]���޾��6�{j#��	;��w�}@�w��A�O�ΜIF&�rx�tԙ��duiV�yz�L��y8$��5Ji��v�:��}}��p	9��b��|�[�I�ǵD.�� ~VI���F�n<rA���/�<Mc�}=�/X$j3���sZ/�뚤V6�o��ߙH�^k�Q����%+��9����V�p�?�fQ��:˝�ƒ��gۚ��Ƹ�Lc󬖺�l��A�����2$�ĝ�O�W3}���[o9�9;����i0��' Q�٘��6$d��� ^�8oU�!�Go���pQ�^���z���� g$F��ݴ��7��wk���4��7\�{2�;����C�5۫[1#;���#�����;���=��JϷ�� 遌V�=�Lz�J�̶� ==�J1�#��D�8�8�I��9=��>�?J�ۿ������O�^ӹ[#����!�TF ��?/��4�g��tso�\�� �Y�E|;c kQ��.y��?h�L�5E]��=ӌ�Ŷ,�U���k��nd>qʞz�q��0�'��PX����HN:�+B�H��H?�C��� �����$�3��S#�=đ���A$a�%��:�އm�� ֩V%�?oqP6x 0���>뀽s�:�1�3��TL���6�f�Y��K)��P���/���T��:��Gz��c`F�9Q��_�T��$�=�18�z��ґ�T��b�L��l����~��>��;$��7n�UFl}�'��l瑙��$��+#�\h�� >A=<� J�od(��J��A�5��o"#m�9��4��S$�'�#�Һ���V<g$�T�I��ô|��:P/ۦ�~�j��
�^Y��bb�O�����g4�h&��w㎕ W��[¦C�wlt��W�|)�����J��w�"����ͻ�~m�E}�>�V:I��dw'�Jʳj%�{�����1o
��>Z�lco\�ҾH�5�x�(���s�k�kƐ��r'��i�|�²�x��� �ɔ\�g۷5�I��kQ�z՜n��i?(l��>�bF�Z"��wՙm}�����B$��j�Cc<u�ӊl�H�D�v�סc���
_F#²����s�Ҳu�l�D�Uxu��i�n'��W$.8oC�Cb�Ga��S�m�{K��.FT�j���Q�b�h�ǒy�U�ʊO1���㩩��E�Ü}i\4$+�,�$��'�k�/]�\��pP	�O� ���Ycn�-�=I�+����ɕ꣎ ����"�Z��]ryⲮ��+��\I#O���Lq�L�O�$�� j�(�o��v�C���b�2���:�ULs��SVUVU�7����i�����1,�r�ܐ1ɫkk۳Ì��eGz�:6���ڣ�P݅�1�0$��8�F�뚨���*�����>�?Zdw;�wsH
���?Z_�W:N��#�nB��}~�6�I��U�[˕$ S�R��qvz��|W�h~�y�f�X��3��>)|X��4�`U
����Wƿ�Υ�x��:I��(��.y�>���?jo�|=�S��=�M
���������vu��;����E�V�X��|��WВx��d ��c�Z�^����ˑ��� �S_@���I��S���J�ݞ�'���3.>���v���q?��ǟX�'���is����g$����Q�����{s�Q9lf�~�iy���?Zw�&�Rgu�c�&�%����?U���H�7ߴo�獶\��p��꽍A{T~���I����7�]��C�1�<��|�"�B�^]N�\��π� �����6�"��½�x�Unk&��#T�z��4��;pQ���7�t��M:�v5K�g����d�V���7�$��>�-��	�_�G��B�3�7g�R�b�,�g��cr��g�5�/|K��'o��>Q�x�#���W[�Ski6���f�2�ܽI��򯛴��E��f�W9,y��TW71��7��oX���jHbI?x�H�/qT����F)D�
���]�9tJZB�B�@1�g�SWlp����<��f��
�zsW4�,�9��)�%����Ĩ�<m�n��X4���Vi3�"��Vk*kDkN���i� �T��!H�>n��h��m�3�^���kS��g��eE�
�7��_�f˔v��1\r�RZ��*q�S��{�흜�	#���^�'�X��as�������{�����`��^_⏃�"���|ؗ�F�*�U��
mh|���?���2&����W6�6��f��[���Ҿ��m�*�>d?��x��vׁ����=+���ʖ�8{Kv��g7��l,ʤ�ݴ�y��ŵ��m������=��n��+{n��Ô��w��s���B�1��j(�¤��P5a0˜3������=i�7*��f�נ�@.7C��w>����H�������S�Ⱦ ~̶��;P�O)X�U���1_4����_jRA��iaϓ+n�O�#����I�H=O�� ��+� Φ�`,�� O�_r��]������� ��uu� �� ϱ8�J��%�瑁��ζ��d��d��9�ދ�Xq�&�)�⢻_2U��$�6�@q�Zӵa��z�����m��X��2:g4�7��=}i�d�MB�V'8���z�Z9���]��]��yǧSӊ������!\s_(x�y�M�#�<���{V��&�bm���=sK�۞:�k�����98�t��Vׯ֜�,ۆ�f*��H�c;�^2 Mp@���_����TBF �\��g�=�;��n:�U]R���Zkb�ʜ�zJ�1��[$���]����ɵI�ST4�V��@-�n�׵z��������sXԩm�>gr;�)b��$U���ڪ*�I��c>��x;�s��,����s:sZ?�/59>H�k{��� �z���c��^ɤ�~�
ǵL�`�8��5 �|��QIlG7��z��{�xN�+���k��W���đ�h�� �Z��X�7ð�#����+�Wܼ~F�`V{�#����:4�B�A�u�e�����I�>����G���BX_�PI8���[�Z?�U�0�L��A�tA��[b=V��+�p��j�q��?�IА�`3���3�? k��SG�>���.�;_�r6�P�\�=� Z�����L�pɎݸ�;���ÃĒGnC�n��W���7�4φ���� X�������|����xs�V��DD�e�~a�����k�S�M�����zΕ{s=ݨ�.~FV]��P�eZܥ�N-��s�ߴ��v��sðFN����~����WX��R��=:�����{7��^"��:�kr� ev �(�d bs� �5�e�I]�`��@���kь���W��S�G��g�.�ᙣ<g�E|��.�|�I�}?«Gk��[nz��Z�r�&��z�4�60�܁���:��?�	�H���1�2?��TrN�
�ңcԱ#��H���M�kS迅ߴ����zL�Y-�!�N�z���� ����"d��[5�t���pR~���L:���X�b��(�SOi#�<}�y<`
J�
r��[�k�3@�K`x퓊�(�+L����ڻ���%��W<�Ρ�F6EFm�M�\,��B�s��\���5������e�k㏈�j�ŭ@���y�_[~�2���v�Eʑ�8��MmOH'����s�5�nF�'�ƳP�k/l
ڷc���˰��y��W�*���1T�_�c�n5ۊ̡�nG� ^��Ҫ�[�ZLT&A����G�|�.|Q~���6p>�����e��PG�W�W�e��E��[�s��k��*6%�h��U4��� ��ǥk_i���R�c����w���˞��6�m�
6󞃠�o�y����6�g$�RGN��ٷG'������4� 6Mcx�b�M��7#��+Z]>�`㞽����\�iW(��7j��Qџ$�2Cyp���;A� i����k��!�"�y6�Gh� �Mx}��=bfwH��Y�NFk�~�OT�t8m�EX�fE>�t�R�5�V;y&*���z����OBO��������Ңo�d�2;v�1�K�,�r���4�����o^�����G����
�� h�Hg���щt��G%�����q��K��YQ�n��W�|Z�?�x�K*"�N[��\��f�_I�R
��TK[�J�wk���78��Zĸ�Y7
��~^��d�� u���"����A�ҧ����ϴmc�����R�v#��]��)��Uw-줎*)>���
�O+�Z\�s/�>��X�b�+���#.��?/���{O�Y<��>p���F?ƪ��ͦFy ֌c�J�j��ִa��kVf��`��ƭF��P��G�N��z�H��B�bF ��W�����׮x��<$mɯ$�iv^���8� ǫc�������c�K��9� 
�?�я�Ȭ2�������E�?����*��B[_h����ֺ�7�4���9����U��3,x;�oֻ/�1��<�ת��}3�º��?^~�/��:����Ϲ���Y
�RH�s\x'E^��_���M
�`:��������XW8�{Uh@##�V�=?:H���K
0��m�[q��OQT���|��x� ��^  �S�c$ױc ����è����u!·c�|l�tu%rw�}
v�8]6
F1�Nּ���G�j�x-a\(�?Ɣ#ʬT��k�e#k`�ڨ4ųۚ����~O��ϸ<�)|��+C;'�I^�\�
���0� �'U�����ץI�������O�Z�����*J��g�ͭ���ݢ)�&b	�<{`W�?��Ǘ�E�و�L� �MXo�66;����ֽ��
W�:Zڡ��<����c��ǎݪ	n��J�$�{? �/�݆H枦g,����H�c�b�I� ���Q����?�Q6>U���/&��5%�@�Tz���
�$ӣ���M�H<W�_� M�ˋP[�E�C����u[k����n�<u5����;�u&=�X�ц��8�jmA����1�z{�/��8P1�+>o��%I,3����,���p��0U�sO��M�ֻS���s���ޫ7»�ؓ�lg�iY��/.�H��y�|#5kN�̿�N*Y�se�4Ԛf�X�s�� _�Q�\�;3�kY7D��!x�h��5����H���jC�'��%��^�)n=�SUx#��N��x�C&8R@���1MC<���+��%��^�k�B\s�����ߏs4uOp�_�H��ƿx��g��}s�BI��;��zs��ҾH���!B��]10f~�s��<�n�I#?SS\�lc���Q3}Ley��␂�
����L��b�c'��
���� ��ɜ񞔜s�2iJz���� �@ǧ�L q���o��� ��S���T2i��ww끊 V���8�WbT�\�w/͸�ٺUwE�h�� Pf�����rHT �@�$�Zl��4ۨ�n���PQ���ہ��J� �9���� ��x��uN3��r���献K�>����.0S����vtF]E������󚳯�����s����Of��Ìs�K�ڑ�w�?Ƌ��[P��o<�B��I.�a���Oo����\�4A�q�Bi��Q����𧲻-63%�EMĜ�s]ڮ<+<w��S��;��G���6w�E��={T�4��|�${p}��U'ʘ^ř�%jP۷�!;�}{W-c,w�w���m,���Ծdw��:�d!�j��cQJp	�����DOR;�-r� 8+��ݕڛ[��Yx���d�H99'�ֶ��7X˲���������@�mc׌��*SO�N��A�a9 ���j�{ʎ�ʶ6�*�\Q5�?? n<� J猟=��sЉ.���gn�/άYٴ�'�9j}&�&��rǩ��>�30 ���;���eK�YY���<����U�G�;��2|���DA_GٲM6�6����'ߊ���rC㋀A�]������U3*'>-W9�8�I�o�# ���"ȹf�y�1�+����K����4���=����x�i��RB��${f���J���p�������Z�� eO�껪�*�p�@����
M=��+���~��xBR��!�M�󻎸�m�7/ҭ]0ہ��j7B���ڻ��pJ�/�n'�8���	��k��Y�>f>�ǽE��]SkK�n��H�}3��Eo��+�B4hK�#�ݏ�_H���w�>���;-�5��n0� }�#񯉾�JO���d���0	�;���>2i?>��7	$�ax��7>�PEG[���>����WM���;eb�)㞿�o���FT��B~��m�4��Y��;f�l@���'�3�u�.���x�H]:����xg��\����r��s�)��rs�{��B�&�S���8�l-ޤ��w�晓"�q��A�cc�E�(H�����Oj^�Ab웲O@?Z�o��$�`��?�� 
��LS�8�@�簬�"��v��^�����������q �=;W�_������1�wK#��0,O=�5�<߹�0�w��_w�>?h�ݎ��^E�H�$`��@�������:)�5��?�֏i�A�{F-U���d�1��&�"�!@��?Z�����f��S�Q��� ާ�ŧ��]���� ��\*��%�a;\�6�9ޣ�����A���Pp*؂�)�����j�!U�1sU�[1��1����W�f�_���U,��;��>�v��#��|/y<���̚L\W��C�X���J��M�~������c��P&ۘ�a�@�V|O�y����3\�du�YY,������U�*��Q�B�zf��}Kc �ɩe�/��v"�Bms����2�nj�ڭu@Rt������bLe��kZ�PV�.j�AfT����|�g�5���x=+�ߋ_5_���3Y���}~�iz�����"x2���so<
��EC�r�+h��oh��zo�!>3�����f��o�׷|J����O�OaiY��8?�ھ��H�RY�qt?J�ݬ�z�I��.�(��8o`zf�����2��O\�a�B�Tt��?S[qƭ������nd+m�1�8�5G\���7`ni�O,�sZ:ncl��Y�7�����@�F~�2���7��?���rG���|�� �_pFBA�A_� �?r�Տ�<v��?�}Ð����5�����#n'�Zu d�Tq���ӦS� �+�&��!W���j�����S@QU>srp*̑����f?l��k@�Hy=i���~X��1����g�y� ���3�y�����n�ھ�:W�>$���V�	�~��q�$Ү�57*��8�ʡ���6���֣�\F8��b"�[8�4�''3p��0���Xg{v++�u���c�4�r�n� Z�ȍNNkJ��6[�5B;_�K���@ �5��p�v��<}3Y�������c�U�i�����6o�gdt���3ÒkQ�/�9bkڴ� ���� ��q^�t�"<|��5�.��-��5��Iݛ��i99� ��5�� �1��5�-�m$�9�ڬ[�T9<S�X�֮��w g���^&�3'*�t=O�uZ�5�m�$ט���%v*�FO���R+s��v�N#?ҹ?X��0U\�U�I&��?�jϾe����8��5�	;�T�F����G�����K�{T���<y!�cp�z֟ٙ��5����YA�1��SHLxf�6��?������3�B�R���އ���,>_��G���&ee�!r�*�4'��i7�c~�`��^� ^+鿂����>�n�K������p}z~��7|Ccj���U��deO��`�~�Y��:#�+��MOFR��n���.>;�L��|�~Ң0�c8�I��6��7`�Z�ٿg}{!ⶔ��A�����_|$��u���f�u�7�N8>�Q�d�5�E&1n�I��dn�r��kZ_����M˅e*rq�E^��-扦ǨݫEh�d?w>�Rp{���y�0�|�$��B�W�|Wo��5��3Ka	��2eT���ះ�^*����)�*��9�5L9���6T�F8ݟ��7s)a�랂�gğ�׈4��BO-Kyq'�qϭp�>�ռ�!Z9QY���Ըٍ4�0 `�YI�x��O�}&��1�W�z�t�,���"rrF0:ջ�{8������Qa�W+�ėv�3�v�l�����ۼ9z��ڭ�?��_���亾F��gv?Z���#{O�&Х�F8?�&�Z+ms�0�ۏs�m��3�X�k�s��{e,���FƜK���.T�׵T��x�j�:�̻����!���UW��J�m�<��Q,|�$R��{�a\�vbG��Ev��Zܸfe pq��m�ǜ�>�1WZm�g�t'� �UWM��F���*����O4�/޳+R���?(���ٰ���~��g����NiDi����r:P�}� ��z��g�Қ��Q����4�ċx��ʊ�l�cP�
�=�*F���RmʟOLS���'�zR�#�~T������+���^�08�Ն%���A����4\�8$�ƿʑm���-N��d�w�?b>� +��m��O[u�zU������!�$�1�y�Y���`�w��X�"�oa;N:UYvy_�m�ptg8�+��g E@����&����X>/�����pk���`�?��m�]�;H@ߨ����MP�����=���$��##�O㱨!�x�U��('Ċ���`d��~�ڐ�3�t�a�eo�xެ�\JGL�R8/0��c��^?�u�_��exb�0�k�_~�O�N��_� <�_�!���r(��'����Y@�^On��� ����i�9��;|Ƹ�ID�q�=��A7������猒{~��ױ���|�J��f���!P��tV�9ɮ�� �_I
r
GԀk��Ly=A�vj�-G� �#�����$��ҬF~c�I �u�ڥ�Q�Tg����O��I���Z`j>
�u�S��C뚴FW֨�6�ǯ5BFe��4�ś{I���S�ϥAbKB}O���WB�<zRH�1 q�N,=8�l��!7ӽ1s�U�)�g֙��� gC���3?7�R�ʞ:R���~����Fv��ҜT:jz��`<f�"e���s����SB��ހ+�gv}=(eNIPj]���"�1�N>��p+�Jǅ�;�*s���S*m_z�5�JB*IwQ��g^BO��ҷd��w����w犴#��In<� $q\�	mr��'$�z_��7 a�\��k��͎~����Eh{��sڵ-�Ǵ�����Ӈ�zV�c2u°>��Ne�R/8�@ g��2l2U��7C^�Z]�ǎ�"��o���^	�q��eS�h%�2~ђ>ݸnY�09�j�6���I��~b����$f��}T�:���!������]123�2H����̣��J|��3P�� ��Tgpe��_֤g�4�p�qɤU�S���bA��ښ�8��RHpH~�ڹ�{��L[�# ��d���}�SY���<�9�by�2��\�*����5i�lR78 U�\��)���"���ߨ�����=j�.��#���s`� p*F{���/��J�Ԍc�$~5�gEbH�[�߉���/�ɢj��`���Ҿ���d�4K;��2F�q�]������B�q�XT�ƥ�!h��ߔ{�X׶�A���#�Ux�c�����%v��x�J���̳n��������	��V��V���s/P:���.%k+������Ғ�C=�M׭!��K�Aҹ�WOqgi��ćn���:�C�|�_n�����sg TU���#��^){:��p6���	��4^E����:g�U�-�P���?JtV-4E��ḯ|F6b,���F?t��=�k���K�,`��r9=1�ޗG����̾Q�999=x��Y�YK��<Y�g�1���Z��~�-ưcV,Mi���� ��f/���9�x>�_���9%��t�<p�?k���';q�\�����/B���(q�s�څV�X�v���g���u⭍�D��q��jilau?(v��u� 
�D���~�<3#E����x��O�m}g�Ȍr���O�{Ƅ��I��m���q^i���qm./��#4hF�y��~��G��b��9E�:������3w9�*_��7�����f2RX��n*��9�idW{�t��6�8��b:�Y[�&rH�9<�՛���[�0���=�*99�#ml�?�Z�=a/��\�O�ցr��P~a�I���$V`��L���oïb�X#bI�O���X���Vvϥ1jlxg�G�������C��y�O�MtC)����Oj�����jc[�/�$��*FAt�E#�8���j>Oؒ�i c�-I���5m�2�� O<~u����+/�!��P�&|�B9��Ν��_
��{y�ݶ<f>�櫖�N��+=�/ �v���/�#��O�߉��Z�Q��I"�$�.r	�\s^��<�xO���֞�������֫��.Z]*7����&Ki��=j���R�
?��yx�^��k���:?�<y4��|�L��Q�F1^9�ٮ��� ��c��t�<�nK6T`~t�%L���yf���]w�8���f�ʍ�6��έc�� Kԟó<iv�#*@�p	铊��ZG�<�A[Zy�.�v����'(O�E>D�g�����R"�,��s���V~��WCT�{iT1��N>��1��B�k,0D��#�z����S�~�O���V� [X��ʑA\l�\f��BRw���M��II���2�����跺�҈S|;I<q�:b�P<'�=�c��y�Ha�%��˺�������j�����/�/�;x��o�2�ʪz{d������ͩ��q�����zzV�yHs�ғě?�&��Kg�n
����I�o$���F@	�+9������⳷�Z�ݻQ@�(� v�Ǿ:W�߱O�㼺�u+�Ԭ-��l����}��ڗw^�E}��"Ⱥ�u2s$�B��?���66�t������E8�F1��sT�͇�hx�XH��>+��ԃ�|��՗�����ē�^��e�-�<��>��%��es�x�hi��v�ӽ L�/>T�9�V�]a���k���r���4�����O\q�s�,5#;�z�t�Cʸ��?w�3ѵ_/n��k��ԁ���(Ac�� l�+�xn=r� {bI���c��_|H�W�Üb��B�NO�~��@���� �{vQ���X�n��s���Q��:�?� �������s���.�BX���t������)#�}O�pZ$��F9du�]���@?)���wC���J�����I��Ҥ�k Ây�����Hd�!g��b�.	�r1��g(u���JZ�c�������_��	<?��s������~����l֪WҾ%� �~�xkXծOc�_p��/��\�gS+�ɔ�G�S\6"#�������*����z2�3�֬��qU<�� ������) 3C.7ߵkIp�l7ȷ�sրQ��ǚ`~1��� ��<����|K��Eu �ϸ�k�J@���s^���"��;[o�?ִ��:�l�^��������l�s��:Tm��?_z�2&e��Sw���U�cׯӚ�䃻�z�E`�/^y��j�*��.@�����5���yx\ /�PšȲh�#�}�[�T\j��H۸u�XZ5ȗKS��q�>�J����e�2_�y�>�ԟ�z���o
�np)��,���`����H�N[�cU?�
�����"�g��dӦi�j��p�pɪ��ߜ��]p�� �y�9��QasZ~�c�p����>T��jZ�ژ3��+:I��8���a�����V�rĕ��T͖9�w�������\L�qI�$m��c^�����8נ��>f$��s^5=Ɏ��\��<�z�#�g񅭶��\N�����'�?*꾆6w�����u�����/J�ɩ:��`p�� 1�����l`�ticWV+1 �{��/���wr�&�Ķ!�-�J����3��s��7�oR��~b��d-�r��Ql,Ϣj�M��>�K��S}�FX8"�O�k����)a4z׈5�5�ă(��8� ����N���=[����IU^�"R��Xۯֹ�ي[CÞ#�~q���M���d^�� �w�6�-�"�]}�1��x����g�Y���2\F�kD�|�w�=�+��'��P�~//��oo|ͺ`G�����]���y�_���L�lJ�Ļ����N=�����GƯ�zV����+�ƛZF� m=���\���o�f�'��CnG�	�_<Ca�����3P�� �#�+��M+�^����ƫO��0 㞘���+ga�&��O�kuFQ�d`��v ��a�i��?��^Oq���W9ʦH�s�~ek��%�� �wi%$�taq��H�s^O�C���~�s��/�i����BN@�h��]nzG��/�?��4��6D
�B�� ��k��H�3�P�l�Q��HT�s��^�w�k�Ү'ҡ�.O�o�.q� ֯�O�H<A�:� ]�fX�i��� }�� �S}[�������ђ����� U]�U��t��|���� ^�iOi�Ƶg�"�ȣi ��@�������R8/������X������0�NH��9�n�W�������H��
�>��������9h�^Q��毽�cп���ȁ��,�<g�?����R����t}kf�8�JǷ��V���3�k&j���'������X>�<`U��sq��e�ǁ�ަ_���*��S����*�d�1��8���ڏߎ�ҵ��y5��e�8�zO`G<�y��OL���&���u���}�9�8�kg��J�QWo8�ni6����ۃ�ӽ+A�Ӱ�kn��4�	���ӊ�-�瀤��/��}�X
L��@ɤU�3�W<��8�ӌ?����ҟ�nx歬aGNi�Z�8��Q��ZF���5���
Ak����*�%�ǡ�i��߀��H��y!z� *`T�3��ҭF��"�m��s�R�a=9�`"���沵��q[sp��Ⱦ?/>��y��a��d-f�Y>0P�kk�*M���#�����瞕vn��U;U�Hl籫�����H-E��Յj�?����Ԏ�!8�s��z�n�A�� �^��!����׎jK��c�~U�����AҾ-��T<R�ꭐs�������H5���|��~���(�H����d,J��`1�Wy�n2�9Һ�'�������)U ��I��M��:Z��&�뒵��?\</��:H�� �x��~L�z����=�-��"\N1Z����ɬ��B�,=G�9��nQ֠��N��U����)���If͏j���T�jL��L��q�Z�wюj�� ��c��LK]�01Vt�+jER֐���3Z�H>ʝ��KR�,{�6����Ӄ�]��"�±[���5�>^�khQ��4��#�{�a*����)��
M��N���t�e!��󊕔r;�(�8$T�{�UR��U��X7Q@�$�zER	8����ހ"��g���V6��"�W��R��*�l��޵R�r	�_P0rj��ʜw�&q>$�F�yņ[\F=��ν'��۹��y֗��FF>Y3\������b���qZP��T,�tJ �� �W�?6�ַ�bX_�u���̀����#�0"�m��W��ݫ`�I����� Rƾt��(]pg8ߏҭ�7~��S�7C-�W>�� �_+Yc� ��
����V����8
�y������@ �f���3������=jy�.���x�*�d�Xt�})�.G#��Ā69��5�o�FA>��1�d���ޙ����o�OL���z��|�1�S@�?��U]��8���T����Dі��@����s�5Nf+�/@q�֬�1����PJ�w��� V�
ı�I��-l�R�#���p6��d��8�����m�V�.��]�<qцO?��K�����Kl����0�}9�}W�ۨ�</f�fH����1_4�B�7J�X(�A�	���ʾ��Ξ�xv���l��<�ҵ��L����d~Z)[#�?ʛ�G͜�c8f�xJv����'�+?P���;�)�A�%WҷНN��þo���$̒/8���ö2��?7?�^��O�٣HcD	�qג�K�jKq��ШH�O?^*u�ԖR;8�������џ옜)ی�������(f��}>�sŚ֟u��D��>n����:w�ɤ������R�p�0��@���?
�%���+�9c���1T�s6S��k��xCZ�Gy|�1㟧�T��<�(�y������k�[�H�>b:��O	x��I��ܽwW-Jr�� ,���$�8 ��r�(�� ��17N溿|@���6���Q^qo:\n�?��pOztb�)���u+���*�zw� ҈�n�K1�Gjˆ镈e}�Z���k˅�[����9�^Gu�xLM�(])*��|���νc����C��:}ݜ ��֬�`���U�^=�Cx�*��P�9�>��}��~�I�͔{^����G\�C����1j�:���ʋ[r���� '���j��,w%T��־�%֓���\ڶ�2�t>�9�9"i8bX� s���d��fY1�P�����O-�����#Y�ῄ��
d�&�Up1�d��!��|�Q�Q�9ls���@��E:#Z%���� ~9�Ͼj�����ۄ+�_��=�/�,˃� �G5�i7�v�	HcԞG�OBNj�@�GNH"���ず��4S�3\+o����`Oβ����۸v���4I�
9�8J�[�	��� ��+"��#0$z�'J����^j�V��Y������������ǽ�{��#3�c�j����>:�����9tH�� ߱��k�u�[��(��	����O�K���4�cŢ�/���Ē�B��� |���5��~	x7Ğ�Q�<���ŕe8P� c��\��Q��\�X�����������)"1�$`�8�� Z�_�R���g�lV�ϊy�;/�P�Y�s�.��/��}�A~��Q��L�x$ 	�N��o��6xkP���{˔��$rH3�ˎ:rC~uFq>�_�+�.��+�u��ghU��a�O\s�_%�ڟm>k�T�r7��/pW�́�}������ڄ^)k�GDgX��.zw�_5x��f��J����eO�ٍRO��rO?�����ZÉ�����W�!m��bF�z�#�^;�ٟ���e�����
���l)����\����ᮗk�����~�W�Z~��м��Z5�wWQ���ab����i�/����+�4� |�Yiv�i[���,d�p=wU�F�����w�g�$�D���2O��b�o���,x~��WΈ�G���� ��I��^
�{�wZ�̒݇�!�_0��������Ԟ��~4҅���R���ec�G�k3<��h�k�����$f`}N��*cJ�NQ*�17ך���1��8r���}j��˝��=)��p�#ހ[��-�֨�D�-}s�I��[�k�1I��� �Z��:�V�0�]آ��_����f�A�g�����?R�A��p[gB@�jt7F�uD1�۷;{�#oy�1`{�&��]���㚆�	/L�{W)e�.��P{�W�'ʌ���M��SO��d\gm6��p��;���"<�W5o �M��jEpeSߊc^�P�<zWM��[�d��ʸ=�zVΓvѨ�$u��I�Sk�����f��?��������x�_XAʳnc�N3���o�<I�~�׳ͷ˳��o�!6�~ek��<Mu!m��1�ɭ����r�A�]��"�s�c�t�Xٛq�������{��3:Ɗ��0h�ȟj�c���Og��!�ɺ0������(����i�H�ہ�<S�폥����k�
��rk-z`j唦9 P�O�R*;����'��3>>H�U��N0��J��	����
��]����3�
�n�l��+�_:Ǵ+ $|��[w�~��j��`ϥE'��t��"o���AR�9�8Ҡ���8>���|c��
�ᕎ��*�O�΢��i��y��ś�	o ��k�� 0�ė{z;�{ޠCB㞕� `���_�,�r��zִ�&��i�N���=��8���۠���x��[���QNV�rI9�j&'�zү|���.{��:9䊍@��z��E�x��4��;Z+[�y�:�U�wpz�5�:]�i�
��#�w�F��R����"��u����7>�d��� �Q���UbI��m$�X2@�})U�c �֡ &k÷ibG�I�$����V(N@������i�#�� � _֪�ʼ7=�̟w�����9�3T3RFA����\K��9c�Z���[��� d/z���.w����c=� ®+RGv���8�^٩t�Jm6�.m�������鲱` �8�� ��`|���VI�w���4�H4��G�1^s�Z=T��;+F���p{VL�Le�4��c�1�ޟP=G�gƭg��k`�yzls�xs�;Vgï�:���I_5�����'�����|IB;��,zk�c�`z�.ұ��Z~�!�g����0���yt������D��΍���zW�/��|�FXׂ��H���B�^���G:ٲ�[�"ߍ<m�x�^�R���,ţV<(��d�FUX^A�l,*����I������f����m�1������=�ц��FV���7j�c!������2������!�A���L�E�,�h=۩�Z��i�w`�x=�5�Kl۠o)�*�#I�2ǲ�T[\d�8��"i�]������G��n$R�V)�h<)�co�N���y�F�sҤ��z�+��S����_�?�B��#� �	��Lc� �k�K�n��K�=�~���2��)նs�t�u�^�Q>��^py�o��2@�ku%��Vݻ^:�9�/�ӎ*� ��j�*v�?�^�$~�%�� ��B��sQ.Cg��w�H�$��q�e�G�	�9�/9��T�s��@������1�����f��! sޤ��z��nc֜�$������x�_ZFb�9"������#�5�0@Z�9nc=�����&�4�U{f�����<+-��cҐ�o'�s� �ޛO<�R���$`�ՙ��M�бJ �i�0 ��'ڔ��CYE�O2�q�Sp5��q�`��?�Q�GZ�*�`�p���=@�[��03�z�|�#N���GBpjXX� ����f,�;���[��5��&=�.�V�T���ms[>?�r�V7��Oj��n�d���k�E���m��Z�����S���[��:Ր]�q�֥e鎕*Uj����P;~!`�2�W��,�d�f��^��|�Ѕ'��xư�����A��� ���ދ����=Fc�R�0�k�)m>A�������k9�Iݞ��S���=JǸ������|ψ�p#��ӮA�~�$s��=�?�{'��n��Nӓ��1��rA�?�v����OS�b���O�+B�+e?g��Ax?�W�'wMa��l\����m��P(-�qS����ڒ���5�wqQy{z�z��/qLl�z�TorsWO��5F�;N)�9}QA�w^jKk�"	ӎ�-�[�s�5R8����k2�kxW��R���c����r=)��(�]�1�Gxvy�l:�Fq�.#FK�i�;SR�U��TUF�c��8�A&��Gn�����P�\gґ�w^h�{���[���ѐ8&���9�����99�[�Y,�s֏�z�\�.q�f���e9�pI5,R���lsT�*�� �V�ln>��>B{�k��3�����3-�+������������$��bk���ɮ �ι��G�=��1ƃ��@ۜsY��|�-Ԍ֌�ж0�*��zS�W���4��⁑\�u�+��.���?>�������p��ۼ@��_��� ���H������g��@q�H� |¿���#��~���i�	�@q�g������Bۉ�#޶�ΐbLg���y�����q�<S~f3�*�#e,6(''���Ƭ����{҅���ޛ#|�z��� �����;SG
9�ѷo�p=)z��q�L���`���M�����=�x�w��@T����q��p0�O�֪M�('�#'���2�8�&ϛ,����@yeU�{�&���7��`���vzz��5�ݸ%�b>���!gcs�]Oϐa�S��#�� ���a��yG�� ͣ�>F<����w9����ʽ��z���l#D1����b����
|Q{�jք,H�D ��~�~��~����Ei�/
���UK���&zlq��|�>���--�B�bJ@=�J���"X���m`=j���+�5p{�]<��ݸWh`�6�v�?�I�2I� ��ڸ�|N���LO�p85���HEA2I�c8��E${}��`*큌s�V���q��׆���$\�<�O��H���C��s ��"�%Os�}*�vK5�G\u�������+�4�?������n�����ǹ��9�I�s3�\��Q~*��09��c�֯��)��������,z�iq���p*��6�q�v�ӹ����[���)�%,s�NM%��뉡B\��A8�ޗ0C�����O�5������x���K�c�	�j�o��̊��}(R%�Լyzж�P�{k�4c�p ���׽|?���#�����o*8��� ���fo����//�����؅X�rX��5�/� �����;�a�o��T��0O<��Vc5�j�#��↵��\����\^K ۞ a�~g��c� }zSf��}F�@+JX��֤i)Gsޯ�V�>��p8ڶ4��[��B������՝mt� ���Tڦ�|���r��%G_^(����6FR�͸1��
�d+�����WA�j����k�̧���KIk;�b�3�Z ����=21Qh��#$\�$�`�`IǮ=��O�*��4�h���wj}I9��d�~:W�a��\����ISӡ�]��-�/kq�0bwB����G.�?���mt ������ ���x�`�n�@xX� 1��������	�_ܰݴ��x#5B2�z��{S����U����E�_�]G�Y�p{t�z�O������޼1c��zT,۳���h6{sJ�[�<Y�R���@r	'q��Y��%�$�9����~*�NЧ���)n �H�q�]n���_J`�G�j���h>�KiFc�v���5�7�B�7ҧ����+x���¯aO@�5���n�0̀>�����.o&2O<���39�={Ԍ�����r>��-������-n5��RG�5������$Z��=�$��a��Mb3t���p��A��]7a{f��n[o�]����i��Y �wV��䴑`��8��$��l��ӛ.��?:�
�'���n$T�9�+)$-�x=s�uZN��k�{쉰T����4��e.��rt��e�ԱʒF�]`z����u�E�4�[�����4}U��v�o�H�8�+�V�O��C]� �?�� <Qk�ZHM�m�炙��� 
�'�j���Z��G׮�.F�:�Ck����s�t��֛�K�t�.�o�@��;����zKY���\r��6�MWq�x�?:�5kB�V�?rw
���7)�\b�b4>�b��^I�#,���4y!T�GN�I�Ef�+^ͣ��z*�1�z��:6�gP�x��Ϗ�9,4�?}���� 
�1ob\���Ƅ��x_N�|����������_8�v��uh�� ����*Es���yq3��ٛ$�u5���������=�1�1�Z���2����m�ˀ�2�3�z�o2;7\��9��|S�;7�pG�?���O>�*��Ԍzg��&�q�ɤ�0��9X� �F�y�G.8�?µ��ڢd���<)�sW���6��6q��j��CLç�nG��_��M��J�H��`�_pFw*���Ҿ%� �{���wU�f'��N?C_k�
��|L�$�J�O�Q̻�たZ�ݜ�Q�a=h[q�D-��ҒH���;����<w��l�MH�c�ޢ�O9��B���ל�^��_�U������W��+�^�@� � �fo��ֵ���ܫ#.��{�F�8�U�-�1�q�i���<���m����Kd�2�������=JڍÒ0}�v?���|?y9_�'��3UdK��� �ޞ��Hrp��,{d�J�'��=��ZF�׊He�Ȏ�#��ZF��{!�|d�`��	�q��� �N����i��Լ7�X&�����9���o#WB8\u�������L���'�]��k�5TϘ1Զ+'O�|ǡ�i�x��}�g�nbn��c\������8��^��^v�Q�Ú�V���,m�5Q�5kk[R�=2=k���,�(
�'�n���䐒H�s��P%̳�j�_�W?�'�5L�Wh\�r{SY�!I>��u���*�,y$�#�wdQ� ��ߊ&`İ�/�)�/�7֖�9�g$zҫ6�G\qQ�Bs��jի�m�#?��E��������%
\^®�f��mT*4m�\���9#:�H�@�PsI����xN���9-�y���A�}6�Ě��B�auܪ9�P}}�t�
Q��31o�g9���*�[�j��YeT8�q������a�kX�[��,1�m�?����t�6����?�=k�XK"���2�6[��np��X�jIJ�.�b֨��O�:������Z�e��v3��㿡���|���G+����}�u+[���1�򟱖e�i��������ef%1��=>R9#ӯ�^�&ܛ8&����B�M>��P��c���RC~5���Q�����F��`v嘑�����,��|��Zw9��)�VP�%��Qd*�gލ���yQ���aQ�ݜ��֘�z{�"c����/�6��	?*���_�Zl{o�� I�����m�5ʞ>\u�� �>��l�)*�lD�0���T�c�VͶ
���cdh[�+��Z� ���Y�ekF<��ء�p;T�p�C�_z���*��ePW��T.7G���"��g5JE�3���@#k�8ɦy�� �Z�.�8��>1��H�� /=E'��ȫ�Y㌊O,�1�@>�|�O�O� Z�ce#pG��=?
s(\�4���$�_���5x(V#�EU��h9a���Ӿ�{���IA��҈��
F��Q�|�֯��џ�JUP{}s�@Q�Ny�H-N�*�8╣
Þy�����<Ӗ=��fL�i�:��y�#=8��T�$�®3|��J��w��@p^,��Z��~�����?�f��C)*0��>b�8��x&���[�N�ю��W�P��p!�� xyWv3��V̞���jUn�֣U�1�'�!5�>��b�gZ%&�����Z2֯�~^�� `.�>b1Yȣ��s���������cp�[8��|O���=�|���0�K�ߚQܞ��i���tP6�� ҽ��Y���&i�!��>��^a���wT\�½��M� ��گ���]ob"~�ƞ\v�:,k���*�<��%��fzlO���t5��ظ�Kc5f,���5Yg���t�Z s|�לw��3���Y��LԖ�n({i��U��� f�>
�tNi6��\��qnBH v��kӹ�WL��*)sЊC2ZԱ�J!W�A�w�E$+ש���(c�4�c$�zg5���4���;�ہQ4-�`J�(0)6S���<�2޴ϲ�Q�iy\d�3�G��R���c8!��Z��������Z��E���9������8�i��^Nv�a�I\����#�j�F:���v��ޚC�h�U�oݑ���T<��J��R: �<P��~��|>7kQ��?:�S������k����g�5�/��;�k�B��hC���P�v��U���f���RX)�֟��M\w�ց��U�־o�ɘ�G���� W�_GȠ�sҾq��"��aQ�Uϕ�j&1�n���_Q�M|�˶3���_B�ԙ���#,��u9_�����O���[����j��.G^8�g<��)��'��Uac� ���rn:T���J���q��|�v�sv��6�S���)G�Fw�*�#b3�'`y<�� '�BNi$��\�:�7PO�jHc���#�R�ۅ�l"��'�Nխ��ve�棼���t��W2�v,ݲFq�4���Y���Z�~|BԾ�\6���J�!�O�s1�ܓ���3V��j[l� �3е?�]Դ���R�E+�wlb��.�ldb�����ɒ�!�
y�MwJQ��������\ۻ�Hp�*��d~��.'$bFS���O�sikQ�I�q�⬯�1;d�=0H�.�畘zU�Wȵ<�����q+�	�ҵ6Ll�2��,P1��2�Fy�HΖK��
}zT���r{o>v�]�북�6�x�Ns���f�x�'<�5����8�/�}jk���|�$� {�jW(Vܹېz���"���;T4��0w������F��L7�'�D���6G8������Ө�����4M����O�+��w�Кa�Q$���������*��85�5�ծך9��=�i�h���	�+Wx��$�
	;=�/��=6K/V���^]c
wc������$���/[Co�x�����E4� ���ڰ���6�|�$N2�N��يA;���z�ѻ��3�c����c%W�+R?���y,�`A����*�тA�ԕa���>�M&yR7V���}�am6牆	݊�e*ĎN)|��LF������Vr9�pz��T�^�5|��e��-ӧ�*O�y�$<�ְ۟�O'��U����##���.�n4�֌����q�A���)�h��c��v>��,�jl�H�
��t�^�����IN� �ߧ_Z�����[�^�o��s���h����5���*ћ�e�v��;��1(��h�h���Ž��V\�I���4v����np�8�j�Y%����p{
�4�Q/����f�A���rf1��=���_z��i?ec$@�~åf$���4R�Q�F�'�n8�� �i=��9=i���PH�b��6 � �s��1�|ԛv��5kO�3;���*�PN�(UMZ�����D��3��j�M]��~c�)��$�����u>�Y��`�<�}i!��W���p;����~}.�]�yyȧ�'I�O��ږ�N9m�y��v���[̻d_�[��U�q���
���7�7�>�kj:^	������kŋ����uj����]���A�j�7�$��*G'�s� ��K�wO��v���|<����%�)�626d��A>�v�f������[L˸C��`��m<��hYޘT�c�z��*OR��=��┚\�w%zg�~��i�n��i����f�B3d����ip�w �q���O��jv>���ͤļH���x�c\��������6p9���=�~ol�iV�.I;�>�h�q�s3��g��c�c��D}����ϛ2�S޺KHmT4mS���V�-�F���p>�"��H���6��F��	�;��̧a�
3�{�]'��Ș�080>�Ui$�J*�ך��ǒ7��'9��� US�9����v>@Hj�3�� ���I��@8z�R��y��q�jR�v_oJ�c���Y~\u5�6,��3��@�u��#�p�5v�� |�An��J�f�R���dN��J��I��Ϻ?`[������w�k�5o��k���5|/��9*G����q���<W��&v2�m匞*	��d�*h��q��HH��[�2��S6��}B;���Rݔ�l(|��@�큱ɪ��3�Z�6�5B�2�;���-I�[>ё����Ia�G��PrL��v�*���?g���ג�C� �-!�T��57G�|>�R�*�����;W���+�7*��f�_ٗFY�Y����ץ}�iR��U�%+&tӤ���2?�T6w� h
�4���Xi76��[&޵�ƞ��N�[(ʭe���أ�ۯ�>=��9��A�;��6l�E9���(�ǎ>�#Z�cݰn����p�1�|7�}	,x�AۧR��\�fw)��~P+�Aocڙ%��FS9����������dR<�p1��ǭV��y�cm�ݛ��_���ڕ�R~�֓� ��џ�U������߳ί��*A�⠛�}�Ӥ,s��� 4[6�5�J�-��c^�W֦��r|�#9�;��sM� ���� Ǽ��+�m�<��E:/X�!�O�Z���?5'����6�3ϡ�I�7Vlb��+��O
X���)Mo	��%�\��ԅ�Q��'��m�h���ny�-sᾳᘚ[�)��
0?Z�G�ºo��L��\��<�k�-lЮ���h$������9=3ޞ�/%r8�'�׻�V����{۫�:3$Lۊ`����~�g3�l�i��8J�UMnrJe��8��W<=3G�	3��,s�Z�&�uG0K"��QN?�W��N�a��AZ��ZFx?�t^�3d(���u�����Ԯ/r�!��rk��M�]����Oi��u�ʯU�޸����vu��}%k�b�HN�vVn�J��m�3�ܕ��3nWnO��S��p��b�s��85&������S���5���φ���ޡ�''H���k�e��$��[H���gӚ񆿐]��lX��]?���Z(؇a�.2+�4�NiI3'\����-��K q��5���?�B��,Ig%�Ԟ�����G�Zy��a��n��@��ӟJ��2;�Jdk���
`[�a� J'�;wg���_�_��F=&��pc�=zc�����6�����H�k�G�?p�L�� ��>�5����z��i�f��V5���8,q�� <~u��#'�\�B4���5e[<
�sӵZV�F��@ˉ�����1.EQ�GSW��l�L��Tsҩʣ<t�rF9���*��F��@�}��$���n85��g� =@¿IDlӊO0�>�Ps��Sן� 1YYHR���&�c�ѩ7�N��y���p�Î�3K�R�ր`V�J{�������2�֔1�('vOJ6��tǥ#a�b��`u�4($�^�}1���J㸫/���*)�=� Uu�9����++z�{U� ��U[�z�L���H ����T���(,2O^z ?�]�%���=S�j��̜`�}M`�#_�z��}j�q��Yv�~���� *�ȫ��nd\��<����s��O��7�����kY	�O�h~�1���^��\n�`8�)���n%=�k7��;�/�g(�9���>.,.l�f���2�����/��߰\	�o�J��V�>��j�' 's��|����M�w)$}Xm?��^�Ɇe>�{W�߲��;u�1"f�Ǩܟ�]�b"~��6�pU@�1��j���5�$����?�X���-��5�l��VU���YB�o�L��H4�ғO8��iy�EeM}���k���'�J�ӗ��U&�ެLp:�i	���#��QɏJ{��C��c�ͤ�8��K�4���h0���(�B�v�ڣ�i`�8��9���1�n��F��h1�ZvߔR6y?�=irZ h^	�)'��}��v�\�3 N ���i�;��ў�� a�i;�ҥu8���_�4��rO^j���2Nj�#iSު�(����q>*M�Fk��|;��'�����%�>X��Ȭ���!�S��s?��|'�C��sڮ9�Vt2�}j�2+u��](Ȳ��`����8����i؁���#��?�w)�8%F܏a_I�1�\���W���7��c����ߡ΁=��?ji���= [I����� C���>�ק�^� �Q2��`���q���~���2+�[��+�&7��I�xZ�Xvh�?�K��\RJ	`B�z�mkQ]5�Vy������aۼs�?Zc�Tq�zZ�s���ӥg큞1��� �Զ�2��X��cژl���x�h����D�We��>��t�c�cP+�`6��^�T;H�US�;r{��R݅ �W��\�	�I$���?L恔.$�&$:��t֌"��29%�&�<�ʭ����m�qҐ�?��1��W���9��k�wZg�H�����R֭��23c�=x����y�xw�DPxn3\B�#A�T1��=s�ڮ"��|��߃���z����m"�Re9i g��澓��_��� ���� 24�vI�0k�� `�f񖪯��''�p*o���猠�H�i5��%�c�C$g#�8�i�N��ğ���h+� �sL��9�q� ���C����|W�����E<*�өң�'u}s�I��|Ĺ��Ky��|�_`+�_�� 	t�i�WAK.��ws��z���ϖ����f���Nׂ:�\ygy$��f�-{�ޏ�o��ך8f�ku�:+�.:�w?�b�x?�LZDC�|��Wh'5�����P��$6��@���H\�v|[�Y\��������#�� U{����h=��cܲ@���]S�O�-_�>!������A���+X��[?�����ÿ|'u�����b0�T�{��.����<'��|L��{f�d$�������G�C���G�(m�FA9W5�5�xo\����Q�q%��</S�׻鷺W�f�n��of�̪} ��S�l)J�����/�� ��a��98]��?�����_	x�O[��V�x���|��A�����x�.��Ѱ7'����5���d�<=v�sInc�e �$c'���U�AK[��3hv�!��w�ʅ�dq�+��_Q|���]�/�7[F�������|M�F]�6��^jQ�2� �$�>��_{�?�ZG�>�X����5��62D�q����ڄ����?j�Z/��/i���ywL����S_W�|;��_��>�����y%%�=��D��ŏ�o���:V���y}{xX�nNG�8� ���ڿn���|+�Y\+�Ҡ
��,g'�~4�݄��=K�� �!�S�~�}�[C�����0���J����<��?g�*��7αښ	dLp����߲� ��~�z����y����$�� ~5�߳>��������\�,�O?�(3���	�;4��o��{�;M���h��!���N����F�i�o�^#��?*%�^8��I �a�~���<!�|�0X�vȪA ��{������_��8�W����4H��G�����lc�
 ��Ӳ���q�)~� ��{�f��Z;�N�Z�1TףwP��I皵a���A�SU��u�9�wޠ�x�Զ���*��-��T��߶�&8���Ѯ�ҀF����ʕ����y�\�|���n2��&��-͑���[:�mȂq���÷LS���l�N�S��Ҧ�<���[���մ����˜�L��Y�63�J�ΓI�#�3�$�5CX��	�� �=j�����s���+{Mգ��Cq��ր0!���^s֥f�V�}$��hF�e���n(a/^���_C֣NW9�+��3H:
��c�zҺV��Cg�&��eWpb
��vVzdz���yWs��g��1X��x��.�%�	xV��.���,5����4����*�ARx��L���=s@z&�+F70����J롒r�Z�"�c7^k�,��N0A�W!�&�:,�����W*���E�܁��̣�h�[�K��鲌v�n�k��y$>8����)��0��$i����x~��J��D�.a�� rA������'��u��j�SHף�-��FRu�+.;�S|�D�a�9����1�nx��Bh�Sӟl��|���ܓ��7��Y�M�����|x$����A�����4����D�;�?*�|a�ɥ����z��ϵ���89�U�$,r2+)7B'?��i�H�G���sR4hBq����C�8'ӊ�&�/�������$����>O5�Iф'=���7����{����K�#J���Ҁb4&��,CqVw�]�n8�I�Ȭx2x�4��b6����vɣu�(��W�֡1���z�9��~�UH*;t��̤RG`��h��/=�>�����<�7|��'� �R�7�g'�<�I�$���{�;� ?˞p�ҵ�xWr�� �>c�Be��E�ۼ�m'��� kR��w�!��rq�4�Џ��o����P�־ʸ]�|���� ���g=0�."�6��W�gd�-�s� ׫�����=��P �v�v��ޑ$2Hcb������l6s��>��$���n�ު݂6�2O5bl3sQJwcۊ �J��o���#Ҽ���ƹ>䐷�T|��y�~�7�K9�	�wb��� e�&�,�����r*�5�)6���6e�7)�����m�J���fx�1xL�2�����V���3#����s�*�w�Ѹ-��V1�z��۳1� w�R%��%��QY�W�6.:����[�ڤ�d,z�e݁������?�>8w��ȩ�����hc��
 jF��Ɠ���J�'��q@����RI	;q��1� eH�GO�J��ܧkg�Ei�g����-�L�v6���5�1��2N3ڦ���)��ƭ�<� H�yy�\��p�9��&ܼ0��Z"���#�z�K0ђE)C�u�-R���$��]
���NrkP�KˀP�/T��C��j;Rh����"��~ξլ�Y-fq�� ��_4Ѯ{׭i�cO�F1��Z�Zhg(��c�>���I�@�m��랕� �����m��x��}��x�v��öC��j�J.�ʚ�?:u�ئ��%H�$"�Ϸ�y��"��"S,v@ٜ{W�]�8;��R�N��pa_z��!QG�׈~����!k)I<��"�k!�H�'�6x���cĞ�5;��џ�����[�G��MCR�k@�ʇ��O^kZx�m#9QV��B&F�$�FsS2�#c�2>�w]�ᛩRx`8ܫ�ֳ���[�{�5�E��q�*��g��0n�w4.Z5f;'���!�t�/��>�����qǰ��^��{R�{���@i�[�'���_�� ���:6D�w�Z��h��m������/<v��I��=p	���~��ᛃ�����+�x���M�/��o*q� � �a�&�䓃Xj�ќ�U/��8<��;iب����U���q�J�k�u�&�,>d�k��?�q[V�y(pppO4���a��q�*��X��:I�/� Z�Ir3�x�!�W��i����D��,�9�(]���w���q�~)~���8��L�}G\��8��B�֜p:����]��^� �^ƅ�ME�#19$��"8f?� I׌R�y�"����8�9�M F�g���gZP�rX~uK���M�W9����U��e��Ƞ<2�j6M���ۻ�R���{Fᚂ�y�֬�\��Md�X�N(��-�X��ڱ-���nS�S��u�ʤqְ.>V�k7�*������U�� HbzV�#h�^�~��R���9�[�������X��4H]@�FB����[�k4��	�5�0�1޸��885)�&R��qϥ|���.�x� �{=.k�����+�a�.�c�?/#� ����2�j|�f��G��1������o���_�t�؉F���q����[=wpN}��i٪6��	g���:�oC�~��?�x��6����o_\�3]\N$l�^_�<@W�n������ 
��ty����0�샯�Օfn9�Юz�{�ȗ=)H#݌k�҇��\f���ÊҎax*�&��~^�ZF��J�ڞю��RK�A�<���up�x�v�Q�nU9�528`2h�D�ԭӓQ!�N,��� i7as�FX)<�����i��Tp��Nր'f���rx�>~��52�[�"�,�n` ��\��2Sٷs� j�ϥ#d�zc������[W 
 �F\u�E"��9��x�����Hr)q��)�?Z�68�z~4��_ҘH�sUfR�N�nF��U���	���a)�J��a[}Q_�*�=M��\܊ZBG=ku)>�H���*["���J����!�����_�0�&�\L��u'45��c�-�����Uv"����eS^�^��ԥ` ~�?��׼,�1��'�E����.<�1���i�6|��Q\n�4���!��5��7���潳��Fm:�1�2�����u�RB�nP����bbe'�Kg���B�{g�E~��sӷ�Q��`�chT8`~�Gjib��}�X2�Z����ߊb��3�s�Ƿ�N������a��0!#�3���L�!�7.02:}}j������u95,�ma��T��m;G�jM������Q07<����ʑ1 � * �������8�O�ȯ���r��a��a�<fxU�����F1�¾J��~Â��d��-�R���O��5+	��M|+�����TK*pP��� ׿�:�k��Z�強.�eo�#�+�l��ܬ��p�W�U��!q%���̬�Ο5��=W�ĝO���~R,�� �s�`���
�G�����]V���Zf d�_}�|�lps���9|�!��fL�@'4��=���_�\>4��I^=�`�`}�H,ޙ�_@�ߴG�~�0o�bIu+�|�ڤ�O'���+ᴇd���I�~�Zۺ��t���#���.�'�����?�j�{./Y�BW<��3�4k_�O�� �:���4jJ�lҰ#���OL�9�0�U���E�&�߉�_މtٞ.�rpGҺMk�G���9,�e�E���<��H�'�.�09�=K>���;����xfo�~���]����H����=YC���\ �z�������9�N�8�=@ռ�}���w4����Ǖ�#�]%��	�c�է� ���g�!\Z�Yc^��z����DC��
LkR׊<�����mN�6� ��Ԝd���5�C\�u4� 1�GC�x�)�6�f�4R�ҙg�_j,	�}(�� �j��i����?���d����֟ � i�>����{V}��~Q��@�������-����|Ð�Sha�E�xRE+�����<|?�zo/l�fWC�9��9��W�?<L�?�����%���� x'�?�d������댜:��m�I6>�����@�\��`y}��&�]A����3L�θ�h�d�K~�q��U� t�������j�sp����fL�Ա� �.ӷ梅L1�Y�:Ԟ$%.��2(���ң�@cC�`v�P�;�4�pO9�F�E=��<���:N�!a��l��&��h��[��s�)�;烚�|7y%��3���-�}d*ۭ̏=�
9���M
k{��.A�ϴ���m�4�:v��ư�I��� �Z�U�1�'�խk�{�0�ǧ~u�k�׺�[ϵ��q�R;�UO�53�ҭ��B�@�	�\϶��$�r� 9��G�޵�]zK�������u��lc����F���i�+��'��ʒ�_5���T�z�K zu?�tW�Ey����`P($Y9�4�h�f'9��3m��}�´m�����f��a�@�>���ω>�c!����ps��c��7_u��Tq7<v��r�:��6�ϸ�|H쬀���)�ɷ���7�߭v^�3�M�[��x�ʹ8W+�q֖H�}�sדN��x��?j2j:�:��c�/j��:Ŷ���c�C��a�Ͻ7��(6�-��x���� x+�5�4��w��S��$��U��6b��3B�eC�1�~��o|a���tn1��/�~"��m�ӵd�v��C� ������_�.�f�;e���x�qG(skc*�� z���kE]'f2G�kM����ÌwNk�TQ� ���Ε����\7a��K	��)q��[���=*E��fp[8
Go|�"�m��N��N�ǧ&�T�:0yҬ/<3�Ol�P
����?G�c?0>��w#��L�C�� 6FX���8ڼ� ?ZϸVVY	�O����-��q�=���6��S�
�;��9��>�]>rѮ~~?¢�5�ۊ��������H�?A�`�+�	�Nqp���G�����'��9�9qps_e�ɻn}��_:��r&����:f�] �3Twnn;R$�0=�Z}�ʽ)���ҥ���� xa��YJ�'�L��̽)�!lq�������VF��zU�e~\�PI&�c�)#��8��W�s�'����Ȩ$��s�Y�? 
*3�)�d`��p=�ʰ��s�U�;29��"��Gj ���k)f��r떻J4�<��;5��_Z.�ڠ�$���K
��VMb�T�b�����-*��:��'ޡ[�vg�Rjb_F��@���\+F)�����-�n�J�����FE-�pp�*��Ts]�᜞Ԁr�
��:6;
��c^�఩��0\�v�C1<D�R�f�\����7OJ�|B�q���镡m��ߚ�f����Y��J�t� �֐�lw�8�1F�&I��n�X���T�pU�}�x���=�H��SִS�G���|�g�_��D��榸���޶�sO��YH�ykqVe>�MV�bf$:��k�>$jVS���t�V���l��Zc��3T�~�:��o��-D� �����H#��Һu�����F�e#�sSL/�c�o;��R]��ş4� Z��
彲k�5��6;_	�kp<�F�HWp�28�} �噉=1��oyqq�C!� �;�N�`O�+��M�>�����]ۙz��zԎ�3�'b��e��	�����~��|����qҽ3�Lʐd����;pN{�J�� �
�<��Ҷ<*#7J\��dg��Ed���:��V��vͪB	������G�W��j!�y
PLH�\���~��P��}+�f�C�7������ν��6����VrZ��v�1ϡ�V�1����V�-��o_z�q�Y�[�2��ެ�l��1Ua�y<Qq0����������d{�}ƨ��������Xz��d�q��+;���ט7n'�Zɻ��[��^e�͐AȮ�%\��8��]W�ǌ��I=}�H>��RI&����	,���{ʹ�(�w��ѩ]:V���|�����KM����,����t�1k�:���	�z��UN~lP��lv�=@���s�QȬ��^r�Z��^��L}��CF�uV 0��
�,�F+��.dY��H	�5O)Ny�h�5?�HH�ڹ�b��lA�?��qvc�c����#�v(�$pjA���k>GҬy���kK
�e?ʪ�JaRsOi8��ިj���~�Zۊ�m���rp{}+���	'\��4���:�������.��N�3����DK�A���U9�8���O����ɭ���=��tb�c��dC�x�Ѐ��T��9�$M��#\g&�� �8BNA'�Ww�rs�\'����8ϭL��|B��bzu�+���z�h�Cmc��� ����r"��r���?���f� �4dq�#�b��g�֛w6�:�VƎ�u��^U�X�-���n9�gں� 
�7WZ�,d"ʬ�=;t����DO���k��KW;X��z���G���Mp��O�:Š��Wi���]ݼ�\�֫���OAV�P9<UXnF����2��֓�b�_��Μ�/�Dn?.:TKq��Vn�u��23�֦Z�6��b�k��I�QU���X�+��n�I7n )��4H��&ᤵGc��%o���i7���RF0y���.�[Ehf�5VC�I<�G� (9��k"���-H5�-@��i�M���9�*z�c^���j8�<�k9]lC�&��!��;��3���-�]��?{�ש-�:f�.�h�w��|��3�?�V\W`�L�]��+�/$
�x�X7Z��o�z�Wo.v���2���lb��WZ�RŹ�S����������J��������[�\���u�w�Mu;���5.yȬ���T�@3��mbI�
y�{ۯ-�H8�<���\�t#����D"��9�,pk��>�O�:�� �G�+��Q2jȧ���=�=ʤ��]�>���Kj��S�­"v�HWy�*Q<T���v�V��9Ҽ�ܞ]�c�_�s_@ {�WϿ�|��{�����h�|{�J�4k��;�<�kƾԯ��TdJ�ڊa��v0*=y?�^?���+�޶��B��)c���=A$��GN;J$a$��u�v���}�MP�bbݸ���XF�����x�g5����k���<*�ޘ�k��[!��6W$�=��b��/5�����5]������/pG\u��)�=�j~Q��ɣ���7��ր��A�҈#�;N���/���$�˷q]�P���q����F+27/�8����R�䰍�'?0?�5��yy۹I�Go� H�0|pO_o��S�q� xg���H7X~��!�d>0�,0ܐ�wN�9Xi\�V��a�!v\}ঢPг��l��/�/��mB��p>U9�5������σ�n�wc0�]Ԁ<*;@��q��Dj��ʤύ�O"�H��MoA��,��0L���q����~~�ռ3g-��!��_�*:��^��c�_��7�T��a��de�[-�r}x����ٟ�k6�
�
���Q�e�Dc�1֓O�K� CjQbWp<~=���?�o�u�6٧(��J�'߭�Q�����C�ǉ�I� j6�I8^rGc��}������-Ž�I8)���pk�o�~�|A���u�a���G_{F�|�瞬�kŴ����o��M�ѳ_�����C�uL@��ב�|��W�'G�?��Ҋ�
��׀H�}���Vsv*Ph�œf�r{W]���f�D7��sۜW�8��k��;����u~@_��z�̄}#�|)�}��
���2=��<:�^��)�&�C��ַ�:�Nմ��4�[�mf�)q77_Ӂ_7k������F,�N}k$�Q��g�\�ֵ�Zї�V��j-���&��0	�W/���l]ۇ-ɮ��dU�\������x~-�Y��������bpy���[�yldc�1��Uo��kZ���D^w`�&��Xm����树s����� �W���.Kk�J�Hb��Jc#��oι���!�������ڪ�2��򫌉��x��2.�
�_�~��m�c��kW�%f
I' ��5򮴓[�$S|�D��Ǹ�s�k�D����쭥+cS�|�EK��6���_���w�\�v+��2Ŕ��J�T�n4-vm;�Z6*8�_jX�ח��#P��4�t�F��d?��xد���z~��(�kl�$� ?C�2�O�5�������U�7Pȑ�^Qa�#pXz�j�E�5�?J������O{�m���M�R>�ہY^.�=�xoI��ۗv�U{N��+Mqp8H�v�O�ѭ�NT|� �+��ױ|=�]���;�h��9�@��^Ya�uk������� t9���:�4���7��7Dg�XǁݪO.������r$F�6��<�c��r�U�5����8�*��"�+?*O�X�.�s�O8�$S�+�R��ψ �a2^�O��+��>�23An�+u�W'��?�?t�7�kWE5��o�p���>�'����A������Oʲ ���os_f����R��3���E��m�������zM~��ן��_�:��_m�3�^NH�ʿ:�e� ���c��"�Y�~f�$<~]�Jr���8�-�H���d�oo�t0M��m�o�����]��A�[?�� %Ѭ��o1���݁��q𲯆dS���:�ԝ,aZ�$������#�T6�G@�#e����f��p����<R���۔����4������O�i����g4���=���q�Q�@�Ҝ�1<q��H�9�G26pON���🍧�X��N�v���Ү|#�X�5����׽w�'��3�:u����`:��)�b��9�_��7�ֈ�O�h��q�F;���񦞾�bh�cڏ"�T�@'�Gz���3xf��;��h��ˋn2��O�J��9��:��F�J��X��l�������~3ҡ��.�-��n$�9�ǮA��w%��~c��A�T<d��TG-���z��:����z	:��L~{�u2y���`�����~5��o��0��{SԾH�C�0~�}:�x��$`�xS��&G�+ml��ڜT� �۞3�4�Þ#��E���tm<n##�f[�:�zU'$��Θl�<�I�B��>���*�q�Wޢ�d�6��J��s��_o�
��O5cO�D'�Rf�����.��x�2E�? ?���g��p+��'ڬ~����ܰǡ����ve�Ё�p��gKܒ�Vh�z�6�������L?Q/� R%����b�۵�棍B�V#`͌�7� #�FY���ޟt���imخ��@(^^�|�7�RCjă�J�u��ZČq��5g*���,zf���h5K�k��J���֔�cQ����ų��N�M��� k����:d���*����z��L�R)Tc�
W��;��Z�o�$��{nw?�EK��<+�_�t���v���s��]�i['޽{�� ���$i�{~�^~�3ǝ�>���j.mLH�6ܬ
\�sR���h��'�)����d(>��w�;���j��Z��9��?�_, q���o�����񎙮#�����Fjρ:��(U`9���=O�-�HV�Ԗ� �q���y��(x�ʬO�5��An� rB:q�9bǴX~�koo`I9�����E�sЌzW��|�h�Ǣ��+��0�"�S�s�c��Ny g#�ط��&�5�>�g�G}�h�G�s޻)<�F�*2��e+g���!�	T7�
���(�(�8���?k2�����v�����f�OU�2�zqQ��9���՗z�[���� �U$u?t���|I�t�KM�@<s�?¹hd�}�kq�������*��c �{W-�/	�;9�\�Uf��W�跏&���<s��_��� ���`X��5=l5�ϛu-jŮd��c,q�EA��F���~�i���j0���#r�Ur�y�q�b��<A�����|p=kՆ�3�U��>�_iJpӦ~�vXC�+��5�zΣ,y72(#���D� ��b�C� ]_�I��ܖ�.�Z1�ж9�W���+A��]j����
��Y
�s��Wċ�_���$����rj����Op�r�Ҷ�G��D�s-� z�',fvq��8���V�;��'�Ѧ��������F��g=�x��s��~V^~S�(�g�=1nzR��:U �v#�*��Xu�0L���v��T*>�^y5�a��>ҹ ��Ih��P��n������� �5�^�op���_��ߴ���� c�J�Hx(�د�->!-�֍��3�� ��JE�X�H��x�na�NEx�|@u�O�O4��X�o�"��/���n�G��>���_ R��'�{W���V�RFl7NkF��K#����v:˻�YIϽb��$l�4�%���:f��L�VPz�PQ�x{RHa���Mt��� |m�ȯ.�����a�qT� �,�92�@��������ц*V�Z�z�ǅWio��MX�Ǆ��`�=R����j����Ve��c�ܬ��� eΥ?��s�� פ-�F�o�g�sg�"Ġ6�z󫋀��(��j̓œ�1|�Aȫ�WPE`�U���C��xzx�uS�3Ϩ������� �R��j�RUn��R`��H�
/�(��9���G� �~������$��?Z��W)j��汤�����ޝs�j�ֵ�|���h�,z�Z�+���S�*�UrO�c�׍M�?�L� ��H�(�a�����S�+����~��w֫�j1Τ+�>��yT����ab}zzR��-�n>w'�}Ec��飑�8�{��6�sUf�-���=��!�90ڣ=h�,u_�`��T��^:�5��,�rd��?�j�}CU��6	&0{V\7�'y`��݇)��Y��W�gi�2W��g$��!��G���l�}jy�c����� - ��_E�B�S�j;4�o�U��kv ���'v;��>\/��x���o����[}ߡ�wծ��s�ʼC��|;���6��P�L���vP�������� ����2x"o��A$��z�������j�a��� �}��{?�bB�s���B���t���ϼ|�-2�A���u&,� *�o�+dʠ�k�/\�>�\���e�7l׸xoőx�K��9�b���T��EԦ��z_��;��K��J�1�5�R��mEWmFx��}�i�Ȳ>�_Z2�`i.|A��D�A�5��Z�.�/#�i�^46�K�M
\ۊǥ\^*�};�X:��#.��s���j� ��
ȡ{�Oq�"�����C�����@=/B��Z�H��9�V�~'�p̢��^�[J��3Jc������E֧Y@���M�4{�x�ܟ��??�&�`0�׈ɭO��{�k�Il>^�暛Tz浩,�Y#�\��ћ �W%���+��I�s��֬i� �V�[H]ZV��=n#R�d�Z���7�^��m�(:zא_\oM�櫺�=��7����$�(�x<��'�vG�x�ݰ��je�����Ͻ|�o㋔��͓�{V�>0�E��=j���{�w�Da`X�EqWW;���I<��Onm�J�V��x�����5?��_����xQXmLL���rW^�n�[�n޵��$:|�$�O�Vڊ��{�z�$��������.>��x�� K��j��&G�ɜ��T��������w�7��B��3��9|{"�<�֯��侇�a���ԼݒNM`Z�ūF��u8k���Y�����=B�Ȑ:���H�a����C�6���Q��د
��C����jӷ���+s�UϨ��f�d\ �� �)d+�� �.�ە�������1�Us.��z� �>Rs^'�|�~�"�9�kb?έ���<yz����s�jԯ��G�ߴ��a�$o�>�Myŉ[P	�k�� i+�e���q�؀ �e9�b��I�ka���9�idcIG(C����RH����Z�E���As���d�egu\�N	��z��`���?1黨�ZO��O�ҙ�eG9��>��j�ôa�)^0�r;S<����R�6�B9���[<��E"<%��^NsN����υ8�����bwB����z@UV9ߞ�;
�)sϦy����[�#��R2�����i��y�2ԑ�E�y��J�b #w'�Z7����=k1XrNph��r}_� Ut~�uǆ�xl�,��ۜ㞣jo��~"��V��������F�=wK��<}c�$���s��W�z+��]��}Ƶy%Ė��$���Lա���6�$:l��!?<W!�'G�<:mྷ���]ʒ��<�+���n-j]����t�a��.a�TG��^���B�s�2���b���bc���^[�o���r�[c�������ω��ͩ�o'��X!�;`�`U�[�ݏ�����P���ֽG���*4Hu	�W�Ԝ��\�Y.�6`���e�[P�|sJ۔���⩤�'S��<��7Q�j�J�T�0G������"�����ѝ���^���i�N�w��H��f���\c�*�[kvmRH`����NhV�G�X|j�]�Ak�M ѱ�����-GĚ�R^L�K����h�����].�� lBH��+;ƞ�|;}��/�$���7�mL��r��֯��Uq��6�r��{�:�nU�����	xj��Z���L��jѴB(���W�0��ۅ}�p��:V����;W��_u=�[��{Pn9lW�5��xР'km!y�4���-c_I_�>>����,v����G-�yRI�T� :ӵ�I�%W�<S`u�2�cr�������\�t� �z{�$f��8�ߜ�#\=��kg���˼,�2��2�x銁��߶���	x���:&�д��n�<�V���tm7ণ}�Y����l���޿5�|Esg�F�7SN��s�zu��~������e����d��%T/#�� :ǑŚZ����.��j�LO237��ֶ�X�*�8�bqV�'�~�M���l�u�q��z����|)��yujn�ym���3].N�|�>k����1e!\s�\W�bx�$�6zw��� h�^�4�|�4�s���|�᝶�#Vgڪ����B���c�I5I4=2�rV�~,M��<[�T�z�~ �f���0���*?
�]b�K;�$�-P���4������潴������G�����Kx��J{31-ܞj��.��H��x��O�fh���\E���]�I�]نc���S�'�p�9�y���n+�}�P�%���F(����$+��X��+j1������\R��I�F$�w�X����naѨOn����F���H-�!F9fS�s���5���!k.w�w�S޿.�^L�9n9?�־���� k+�ƥei����0�Q\�)�Ƒ���b~���_	uD��0p�OU�������X֜�e� �' z�z7��Vxc��^�sķ@32�@�:W�� �O��o������,"L�����ք}�
MX��tH��}�M�!�H=�ɜ/ʼ�͏�#s��WQ�I|B����:�Q�;�?%]xV�#�?�r�yO�G��#�jd�9��`z�3g<���lv�=��R��8�j
44?�ު��<O���Q�4�,m��	p��K�ɶj��QH�.Q�R�ќ���wyaG'��빎
F;�ߵP6z��� ��'xi<�G�q��՟�G�5��-cy��(�.���<W�y+�V+�sV��D�bv�w�z�`��hy� ��v�3����b=���I����4v?1�Oj����Q��?�?�Hx���2���M��G�1���x�C����63�}h��2� d��g9ǧ�Q[1� ��.0iw�w'���Hُ+�=i��q��ҡ�J3a���?ށ2Nt�w�zq�i��`	*�Gc�jM�Xc؊��^*U��#$t�ݞ�� ^��dŋ�j�a��x�����j���c���U�MѰ���}BjYq����ȭ�9�n������Z8�u�5�w�>�!*���5�I��IC���p���{�	=�!P3J�r����!>1��ڝn�qim�t�L��Ҁ%}��H���i�� 3�&�yj�t��/�G�`��.�� >@��<�\�׈�(�*��#��v1�U�z7.�N�>�H���?��F��|�x��^c���k��4�q�};�A�W����#��4Q��=q\ŭ����]�,�����Ơ}'�~qҤ��i���a�LڛF�f�¥	l�K;60	4��۳d��B�ړ�-MD�v�&�4.�ǵ!���ګ�չ�PG��0�q�ҭ��&�-P�y���-@І�����Ǹ��M�E��Q����V'�W�=ϓOQX��m���z�'��&��9�Jt�d>gL~"Fw�@X���l����xf��O��*��r���Gܧ=Fq��eI<+g$�0������H��V�j>R6�+E�o�g|�n d�����y�n��s���� 
��e'�Oƻ?����֪��$<�}Mr��ټ܀?�������{4S��'��X� ���#�~M��߃�U����3��v9�?F�~� 8a����oD~q|F��q�26�}�s|��cϦk{�R��L���3'�8ι�èU�9��8|(���2��Z0I�O�1���"�@S��O4�Q�3�ЂU�WnO��Z�HQ��LU��cۂ}3Y���m���@��s�ߊ�z�E��(��9�a�0��m�*��u�W?w� @ }�>:�ȇp�j�2���%�NgI�`����,�1����/1�#>�#���m��� �@��&�����tl�=���~=M�����$��wm�2*�����4���1I��t��jV?B4/X떫43��3�_�Z܎� �c���� 5/^$aȷS�wp �j�o�?�|Ab�<ʲc��g(��{'���ʜ`TM�20�}9�y�4�v!�b��[Θ���|�Z�2=6Mm�� �U{��̪$�k����&H�8{8�74��}��7tO�e]���o�X��%��'��ֳ��5���h�P/\��y������K}��A��������X�I!�\.������}�-��/'���Ҵ��x�n�U�z����>#[�*���w8�j������VhYH�8ڼ��\S�t�8|���x�I-v���=q�VG��Kc��F��"V8]��������V�:3����;wg}4$��^9�.�x��`&�������o_b+�-|s%�7a��U,y�*��K�k��2�o� �\t�*Y�gF���������=�M��k�Q�o'ש��ƾ�.��5��:-�����$x�0##���Ꮚ.b�e�|Q.K� \�6���בbv��eG�ɭ� 7����x�N����(s�J�	�(i�$h_Қ�bv=V��h�$�F��ix�Ć8e�L-Hn��+Ĭ�Y��!�2���3T�OMu�g�ܮI�ԣѣ��,�� u&��|T�<K"Z	���+�}9��t;ȯ/�H��B��&����:��Zk�S�/<��h,}{$��`�>�bjַL��O���? �Z}R�`�rfP	��ދ��N�u'��m眶>^�)�#���.`���n�f�<∟L�m�#��n�9�8��$Y���[�r$S�O?ʹ�x��*��
�dc���=�L�O� c�J7���~\zԚO��h��FV�ӵ|����I2X�O�^��2�X�[|�2�vJxۅ鏠?��M�@x�V�#�㸆X�c��G<�Hڕ��c�/L��C���lV��F&�@���1��^��R}/�r��ʲ��UV팚9�-�K�Ķ{H�a�5��YI�;r�W����a$i��N|ߴj�!\���ؗ+h}LڢK�)ld�^a�/��%���X��5��� I9?Z��|yMgC���ݙJ�pz�Z����q�(8*;��_m|�^��/���$qѰCҾ)�S喐2��n:��g�_��ׅ��4�,��ڝXs�B2������������ u�=�[�߼O `�ּ�W�ˏ�ϧ��g��1�#����?�E���^�#�$0��lr��z׊x�a��,�n��,	d��ֲ�MlT����o�Z�[��J�?�����m��H��5�N��W�Җع� |�U3|l�YY�� ��U�1sa>��\Ϲ�2���{b�Q�&���k�JV�ݬv�H�B�8�Q��W2>��/�|�ϵu�x�|g�Ƥm�#�oƾV���S�Z�o�y��i5��j���������>c�$����o�̱�ع$��</�j��ői�2����W�xGX����#*>N3�*Eq� c�t� G+y�in;���/s�������dc�\�#�Uۿ�^x���Z�m�bR9"I"�����Z��� 㫏�c��p�YGE�r ���N"��F�g�v�6q֮�ď�x����G �OJ��M��u�jVН�$p7�J�_I6���n[��Y}��TI4�3�<k�5��I�/�Nzב���I�Kۦ�dl�� ɮ*�Ǘ:�_1��j��<�VЖ$���ߎ��=O��wPɸ7\�Q�-�b�b�j�_�&��ov�6RB����e׼]�ukV]�+�x� ��*�J/���6Փ����][��61�׋�|lEs��=i��ZS��9�� �7��6�>����$�>٦�B�s� ����<M㧴��ۆO�Z�y�l��;2O��Q�j�]3NNM�tՏp�g�x��h��Y8�_���C�V���q_/�Z>ַ����� `׭�#֮��f�AʦI뎕(��u:����s�fîN��q
=��|A���U��Yd��8�Y��U��ʩ�G<�Y�x�F�ǑGwr"Hm�p}>��j�k��~�P��S_+�2��ס���fJ��_|R:�8�O��=��Y��;��������g��Y�ֵ�[�7�=�|���Z����>\�<`�t�^�񕯙h� ��ZV@�{욕�k�W�4C�Y"��s^[o���n��˶�ݧy8� �=x���ϙpJN�<����9��>�Ե{U��$_�5�>���Ǹn���|ri��m�޺O�\���%����y��6�YE�l�?�^f��j1��5�|w���X�j���~��K^su3GQ�^>�����W]Jk/�zUm��f8f<�H�<����J����b�3�kd0'����؏zpe�m݉�M9݃�=(��8Ա< ���E�ȭ�@W���/]Z[j���lc��zOj����4����g `d㏥ 2�#L�����֮�O����O�g��n̓�Gj��Hd��+�26� ���\`��� y%��z�c_�\�g8�zR�7��� g�����zŁ��н�� ������c�YG�B�mVB7'��09����q����~���-��%��d�8� =+�@"�hۀ9�l�;��� u�K\��OS�O��7�Z�b6sy� 70۟�|}�Ux���'��k8�q�K�x��ysGs�̢p��pN+GT� ���{��}�(��)��|����	�[���Ҙ�� ���?j�ğm�-�C���˸��{������Z�}�'r��/��[q���Q�rO%���"���n�7��j�%��0��r��}�߉� �`��YL}���J����\�2�I��*x9��x�K�=��WBN��o�W�/k^��O��hY2��ʚ���ƹ���&���#�N��'��q�-�4e��2O��T�,���-ޟ-.],>c�;�ߴg��%b6NGz�ӷ��_�о<��ċ�F�?.�?�B���� ��O.{eU�ۮ
��i�����6�|-+7Q�Sj.�硈�.ͤ���@���c�ػ��'�ɮ�M��|Gqn^H�&ے���ߜ{�_��	��w���{n7��b?Z�KA�≮�P�d�#V�[���?�-4_J����P���ҷ|}�6�ט�`˃�k�[X�|]�����M(!�������5����YFG�5���_+8Ƿ�U_x~����lo2i9-�5��ԍ +�� ��U���~��%�E9� u�q��ٷ�t��?�7��}���_�t������GN��/�Z׆�E�$lq���Vo[�Z��Ϙ@�b����7�:]�6� !C� dg�T�qs(�x�nooZ�i�c�wqZZ?�h?��x�@��ڢ�h�#��QE����{
V(�d����Z[�y#��t�t�J��͙�o�'>⚷EX)�
�qm/��I���$��*�2GL�/"0�v?u��Tv�'q�4^J�Uz�y��_�fu�~\%Fz�֪�S��G	��v��o��y��W|q��Lq�S��/��r����U#�uV8��|��+��1[!���y�ǌ����H�����i���x��}�©�}jl>k�%vY(�Y�%Ċ��W��9�X���V��r��>H�@��Pq����k���=�����$�5b����GL�)�4�^mH���®Y�Lo��1x��V�7?�^��Y����3��
q�{�ھ��w���F�qkC�2��s�p�܉N����fη�I�������Z�� 9Fޣ�������.��vɧ�����?Z��b���d��rq��Sԫ�v�Y���53.� q�U�Wia���5;Hz��z,�uHTrI���Q�Nz��f�� �"�H�ҏ+�1��O=z~��w*�o5ꄶF��P�����v��3��1���k�^��E:�� .���_xf����}`��4	�+.q��j����q��if�$���z���\./dv���玴�x�e�`T��[�Y�?w�9��A�z�R�c[�����p3ֹX����c��:V� ������c�?J�U��y��p���)��$��!�@zT��W�6���Mc.��Gi���4ۍ.��~6�b�X؉����xw�X|)�^"���;���u_�w�#�W��!����)�	�8�+�[ɴ?źo���Q>#2H���Fq��)���H����u-o������#�����ʮA������zw��"=6�%���2pG�A� ����k�P�G�+��A��4=Ɍ�����y��t*� (+�Brj(~f�H����R�f�
��O��JE�� �p�)��֚���=��[��>�|R� �GE'ޮZ�d������z��e�=������8)�~B�q���+�a��0Eӓ���wW�v��w-!9b���`_���>�[�7{�W��	R�Gj����{�c�,g����8��w��
n�� Z��FU$b���u��1�g�=�C�hվ��R�/��&���-ԍ�(��n|7i$�lJ*�?Nu��CǥlM�X���UL��+�g�E��r�Hf�$Um���2x1'��$�+�?�U������1a�6�x51��=����<�ꥸ�7�HF	��n*~$ y�����U��gUaߊn�bH������{���@�6����m�rNjך`r>�����W'=h�� ���R�|d���@�!##5&��@<P�\��9402�F�f=����@/�р�����Yl�Ks�ڲ����O���P�7�ێ�����<c��B���ۊ��ǝQ��ϓ�g��zW��]b�m&$���:qP�_a��KyL|���)8�"�}1�;@88{�Y/��F�:#ܑ�+?Z�4����o~�� �W���z��sm�$��۲3�ǵ\)șMZ�ƿ�*��ǜ.1�����g t� "�?i���+������B�?�sQ�� bYwt���f�����.[�ӷ;���Ɯ�m�V����'���_�3I>�D�s�s��S���E�6K`� ��ք� "���&�ͺX�	���<Qp3�r�s�֘�6q�^����vV�Q�3ޜ�gq#��拤?7�y������PI �N1O��X�-��u�����w9�Qp*pT�=�*P����?�˒<�BL
X�\��ǡ���{8�����$�A�>�0�\P������0&%��7t��*Ο�����ȭ�l��P���H����b�qK�f����6�?{�jxu+�$v�1�����"�|�\��� 
}��F�n��S[�F�i��錞O�v�L�:�Ipe2��������]�w��
v/�-����y��Φ���m��W%�M���co=3Y^��/"�݌��W��#�����3��<`���^�u� 
�<i4��v4i��zWevu4m�P���&����ē�O�_�e�]�|���c�� =?¼��X��_��#���3���U���O[�h�V�e܅��=	��V�I�����R����h�.9#��B1^�j�_h�Zfu���W�~Ԛ��-m�[c�O0�@�ʾz�����s�lִ�F3џN��]k��ܨq��� \� �9�)���G�Q��iaȮ���+u�m2��Y��:Ԟ8�yuky-����d�G�k�����mง�w/��{W}��K��k�/�k[<��mm�{�� J��  �7{�71�������]���9���ƒ�����C.�rO~:�ʢZ��#���mk��7ѐ�,ŕ��a�s�R1_#.$�%i��NT��J�+�׍"��2,-KfF�d���?O�_5�w��_���º�#�g�|E������	9<qK�8?��Q=��8/��?��៊���27 �d��z׉���M �����?���FM)&�\u���,��Q2r����&�������<��Y$y#7(�^�����=
���܏ƿ@>���ڷ�����ں�����3�l���s�m5b��ǄlZ��ҡS�;⼛���.��L*�%W���Z�g�ƕ�5�i�|�H��h�^=}I��u�^m{W��w�,�q�u�%r*h�=��U�<bc��v���I9ۓ�}?���L��<&?�幆<�\�p��_8��o�#-��To
{�xo�������A8+$3 �r9�K�\��c�MI
���z��u���Ι����ۚ<A���K��E�X����t�'�u��TM'�Î�^�AZ����.�l��� h�>P�����b;�|+=��+[��X`ccs�J��i� ��y��L$j�p�9���,}��=�u[��&}��D��'��	Y+�8Z�nT$-�U<���
���6���OO��m�,0���I�SZH�D��T�Ƿj�G3z��W\���{TLV>��0y���I��z���1
 �皭Q��H�
K(�N=������|U�;[����I����H�?
�/P�UP�r���}z}k�O��4��<o
��ܹ�k���Q�J���7~��?�~�kV�$ڦ�$r=��|Mx̳�Q�F9c�����/����<u�NUm�	)��s�|����!�Ȁ|�xUa���x�ؤ	Y�W!�7t�[���u�w蜜�}+"�f�<.9=:������������S0�0Z�o.6g��\T�f�qlu4.�,��Pa�j4��&��,m/��ry�|���lf�v�%�Qoq0�ط�}��_<|���$20U�u>��l�ۿ�:/�������5��mKC����� ���o<%dn�-J��ܗc�>��~�
~�c��%���.T�Y�h�񍾵_�ީ�������?-����w���!�M|�/�uM/�-������w#ƪx �1���c�!���?���+e��kX�1�sj� �: �g��'�?k\Z诸s!��0	��{�w㟉|A�����Kq"���H,p{c�y7�[��OxzR�f����$Z�wFr��k9��x������� ^���� 	��#��$q0>�j��z=����������_��e$�x9��Z���mla���o��io�>��2q�w���G����ǐ+���8�[�o�[M;VMkJ8�F�6�p{� :�<U��4뇒m�g�=A'�VW-�l|�u�+������3��S������?�x����lΌy#���k��|:��-���ii:��F_q�t��&��xOG����쩪D�i?��J����Z������[��Ͽ���_��ᮓ��D}rV��O#��q[�	�� ����ۖG���Z��L��]�����O՝5���E����U�D�-D�,]$s�O$z�+�]*�Cբ-�5�s[zǄu�.��X[o�=~��~η1����k���!� ��s� ׯp��m�~"�=GkHc�<�ʪ����|VO�:��� �wQih��<3(�����ӽJ�7>7�����I������Ÿ�NI$z�k��%0Լ@"�}�a+�O9 c�'�/�ԟZ�.�fb�,��9��=�W����k_��F!����[D��=�⟂� ��nUp�5q0�NK�(��Fb��E}%>�o�C�1��]�F>a������,���'ݸ�����̍=
W��4_&��,��~b�׭eh�lo[�3:~��{��>���ėZ��������v�V ��^j��O�uk�u���|��cnOA���绰2��,���ϑ�+W/��^k⨭f�± ���BG򯥾6|b�|tm=VK�Eă�"�1�����"���Zꦯ����'gopjE�x�<r���� ��Xg�H���܆�l�Dk�\Hػ��,zS/c/��g�X���o7�i�C:N3�6�إ��N��d^��-ɤlm���h$�w�J���O���3�v�e���F9��b�>O'��ǎxv��<�K����=�`m���Z����i�ҀB��O�b���#֬�p�^Σz�h�դ��=�˼�Ê���F�7����aW�⚡��d�ƀ.�sY��ێF{Z���yc�����Y$2G�~l��[Z񷅉�A'��(�i�Rv��x8���EuܻG�=+f�R�a #ޡ�K6��٠
���x�7a������T�k;�L�n�ֵ����Lu���j��ɜ��Z�]���)�χsjڂ�ӄ2fA� Pp�s]o������jV�mev��e� �|@�+��s}����Ғ��v�<��A����r�gɭ�]��ֺ���j�KE�Ok��Q��X��ֳ���Rڞv`p?�gC<���N�I��eP��T���%���E��4��]$�a7s�֢�$^2i#���[ ���*�Kˢ�)
�g־����A�W�n5Kҭv��(a�3�|��I��y��l���cK�1�rq���O��7�T\_k׫v�l��<�۷<g�yw��$]K�=[Q��q�W��r�`י@�j�C����>�j獉c�y�i=wg\���ў������=&�6�. aXg��4��y��}��9☄�W�#�k�����tF����Kq�Zi���8o^1O��X�`�1����{
[n{֝��c�e�H��9�f=�=��x�7q�����GE�?Z��MTm��Ӛ���>мa�'���숎���[P�ݹd��҇^���)+n�5i�M�t�'�m�H�hp�#��{��6a˫1�ι��J/0�n?��2jZ��;���ϧ�(��.��;V��Zu��`�5����ee%O���v\����9���������^�V�G��;O+�X�����,q��Jc33�O#4�s�ٟ�o�tY-��Agg9>�8�Mq�>�o�x�_i7^\�N���?��d��X�h���EF�Ҵ�i%i_��["Ȇ���M)27;���K��9�S��K$μ�y��9�z�d7Z�J�}kSE���G=G�d����� S㺖��s�P2���$�����"��D[���N�����#��V~�4l��4��xOG��w���m"m̙8l�J�~:|j��ˣhLm��7h��#� ���'�`VB��Fj8�s��=y�N�]I��J��H�x����ف���:r*�ڙF�Կl}��͌f�R�b�[�z��So<>�,$�Iϭ;�&<n'���t�v�|��gF�����q[:Ǉ�d�~A$	�q��`����?Ƴ��q$l�h=hb�E���ݶE��3�{���"���^Y��Q�n��3�ۧ�k�h�F�[�zI.dy���5D5�n���a�*��0=����7?1�5�������Z�q|�MǑ���ZL�/Ȃ2�P:�c��u9.H���9����2�y� ?����x�	����iӎ���R��xǱ���o�\�̭�6Ns���d�q���wI$���� z���Z��Vڋ�e�����U���'�ɬ��vIe�B62@ c8��bVq�܎��#�N�bf$q��4�=ϣ>,|_�����i�3y��r{�q�^Y-���
���c�����]E
��S�����_�e��4���m![���}�v�|��'��O֭��X,{���\����H	P	�}��[�.6���p��>S���O��i_��ں[]�hX��0��ˤc坬���N5�X�O$q�6��zq@�c��j�, 2銋O!��9�����[�V;�����O�~^��t~�~���䭜��d�*?ƾ�h�1�+��"C��K��u^������<�Щ��:z��1lv8�ڰ,�i�/�OL���U�Z@h���ⳛ1�$�ؤ*�2=��u�L��@D[p'�jd�|̷9��Ni�����2�ڀ>i���6�ք��!an�q�@z��f7c�^3=2��)��Fcn`�Ra����V&ǖ3�j@�<S�<c�{��wA�FUr4 ��)U�_����v��5p��^� ��1>��N��r8�b��G�?��.M G��g��8�s�欶[�OZ��]�ݞh��q�� Ա�,9�H�ޟZ�ns�~J�5<c�ޘ���s�I��,��.9�9�+�i$�F6�ɨ��Q�M}�F���[YR����Iʏ�l����cs�q��ǃ��xu	V<n� ��?3@����~��[x�G���p�e+!?���,���ɵ��l��x��@�+�>0h1�x�H�f���Q�?J����B�,��<1ɭc���n|T���2m��;��k�&�}Υq#U3�["��g�2�K�c�Nx���&�u��,�d�HR�i遜WM9>�畯����3�����F9��T־�}�\I	N�J� J�_�����̈d)�㑑���:����T�����b9 xGÿ��x��{YTD����q�z�]S�v�E�t�=�c��{Wֿ�+�<mV̫ŋ A���?*��ċo�-B���+
 裑���̭`�WS�ɾ�\q����D�c�r?�� ^�{RIU���z��P���Ď1��E�a���?�����7O'Ɂ�Rd������^����Z�~>^3��}���Oo=͕ԟ+ŵ�1�ֻ�>U�4��X��#nrj'|�c��9����Ԥ�7�"u��*�������9�0+�/�.o�D�LHS\�2�g���F�������!%���j)Y�x9f㿭�Ty�������D��4�6�9��5�~1�as�F�kI���q�}_��C�:����%2r1�\/�%Y�h㭼��b�FN��|�o"�*���`��C�c�3�U8շ�n�Z����z�]'0��n���iM�9�G�;��'z�bT��S�b�����$�3m�3�R������� �P�͵�8<�q]��uķ���#f���8����U��x�jͼ���:��׌�z��ϰ���c�C�3�q�Z_�ZU�ed�~���~��������/�^N<���r�:}���$�6�q1���s�j�~(I�Ȥ\0��J�����h�Ԯ`����z�c�����H|ebn"�Wjؑ�3�~���έ�Ts�Vd�/>�Ж-��n��"��e����cTs�ݖt�Zm&�̍����׼x3�j�h�\�a�� �����I=})"f����x�()n���.�&i���#$q���{�$Zl�q�&�ѻ+���c�y]]2�%lv��WX�_�BĞAc��Tb����|]�o�K4�Kvo��F��:��`ZF����N�LD��W�=�N�Fq����o�o#'��c��j��E���s��WS�_M��	$,�J�a���T<E��~ -���h��~s�|��5�x�\�ֵ]bx���{$���#1���Q%r��=���:m峖��q�}Ƕ+�R�,#��{h�Ks���^��!�0�v��S.fP]��׵O�]M=�=�_$�4���&!f� _9$���^�o�w�z�~���N@-�;�G��(2�pG�\b�d��$�F��%���?-}�o��]�iz���I/���I�#(e����?+zz��*EFN'�sk����ͼ�Hg�^��6��CPX���ӑ�����kZ��S�y z���<q���̋+ue+%N̿hw�8Փ�7֭oy���^g��=k�5�Z��7�qs'���N�s��e�����q+M!������9 ~��V��ɱ��Py��Tt�[��j�x�*����ѻ�$U�L�O��8�׏� W�J�N��j%a���y�*���'mE�H��f1��5���� ���?���}�G��� 믏��c>�c<{W�|7����=���k"d� �;�=X��zR�>����6{jڊ�G�ȧ�
Oj�Bk��3?�P9�'󯧵OڃX���I�+���"�hې��w�־r�ƃ'�5x��M��k�Q�)5'��b�Ӟ�%��L�*p�r0:�@�ˎ��30<��j�2.�]=әI�� *�fs�Nq��������Tm9=� *@t�Կ�u�;�Ns���~��𶣆�R9�69;��c�ix�!��F��TN<���Q*j[�r�Aj�.]fey�g���׊ƛT�����o�FK���������T��p%l��s�z�{��>q�<s�J��\�^k��S۽��kE�X�����;{�ip��4s�C��ps^I����6q��Q4�̪���*��1=qV��r��W��ӎ��=j揫͢�,��Nw) u�}�o���=F�u��3����៏���v�o�W��؛���I��3�_9:�ų�rM8R�Z�Tk��>�����Ӌ��׋n|��A� Z���+�~.|V�~3��MU�[�)Ȋ ą��'�9�6Ev�I�g'�ztq�R�g?�4�!��h���8����%��L� �bŸ�O�zg��T#�<���e!��KV=:���ҽO��>������ǖ>c�Q�d~��8���gж� I�K{Y��8o-��?
�&|d���c���_O�"a$���2�o`pq�y{ڍ��'��V,��(�\�a�X�U�F9>��7AԐ~l�}*�V(�ֵ�?����#�v�Y���Г���n>ce{/�O#w�{W�sx��>*�䑤@
�pۻv����wL��u8������5(a��vQ�|�@�sʒ������4� �z?��3�Zّm���E���ʼ[�_��$-,�r˜19&�q乹b�L��&��CI�b3�֜i�����z�����wg��� �:�>�&� ���댜sۊV��n���ť�q��}*���m
q��5��bO'֟���4�h� id}�L�T��]�R�Q�+'.3�d��
�(��A<d{��Yf��5�����w��=~��y$̫��S����jnЧ��V���$� �U.$ۻ) ��rH��i$7 ���ǯC���q�n�d�zq@��?�'y`��晿�qDc�� �PǐH�)`J��#�q�&�ǚ?� .��p=;���'��Z�byӭi��1,$�2Ҿ� t�Λo�`|�3Y�m �zU�&B�NO>���5�g;��:dv���I�\��֮�hd-�r�doސ!m������1Hړ�
X�8��Y�YTu���N71��ǽ+�њ�)qڴ��i�f����|�?�t:Pj�vy����D�Gl� h��m��%�G�?J��fK�$���4�^����c�c}��8=:b�����+�ԡ�ۇ�LD���`�z��I���x�;����w�F;�d����dT�f��{[�=*k{�4��W�J���g=M[Ҥ���듑LF�ە��z�Y���^���m��ʏ��JX� ����{3*��G���I4S8�+��$Y-�m�U�9�[�t�����|��$��c/���޸�ҳ���4��q���juo�p����=?
���~$�� �M����\׍y�X�ݟAR��Im8h��g�U�ohR\j�]@���3�<W4ѼO�}k�������<�˂OҹVݽ�9�LF��٤۞�_�rY�e[+���4i2��G�O�L���x���ҝ�]��."`�w/�<��0����gݟ����U�	!Q�G�GR}��w��C��,*A�������8�Қ6	�4\�>spw1�W[�Ȭ�22pOӵi0�>��7p\���+	���*������Wa����x�a]7WOc�;� ���x�71�Q۸�g&���de@�q��Reu'���Zd��:��OqQ�YKd8��g�W�����M�v����y<���ە1�޹�p�p*��a�N���g�4�� �߭'�vd-��G'֘���ɕ8�t�y����ojA��
��3\�<b�C�}����H�2I�<t����,�P�_���v$�u���'��RKd�����n�k\��Q�n���].�����P���� j\�0ߕGш'�i�~\�'֘/"���g��$������;���x����o���@"�����w�>�����*O�J0�Nz�zҺ�ɲ�����s���Y�Gn��~��ԟr噽��:���*o}���rKs��l�� ��.���@9��@�@��©�==�z�	"� %� �w��՛1��p8Z�4�uX��� �Ɲ�)kjVU�<`���J�ak�Ny3�Gz��5��
�U�̫���麂Ǣ����<�����ď�`�̟��n6��J���� ~���� ����Zs�����ؾ_ʇ��~U��:����B��jj��36��Ҡ�sڐ#(6zS#�'��3ev�)��d zP���<����n^��*k�y`��Q`v��h���̝���cM������}�I���NuV��S�+�jf�2)�р��a����) ��m�9?֡�H�_ʥ��P ���1�\s�@c���+.�`���c֚��3ހ\'��)C�8Sw�q�|����@�>z��=*�Pd㩩ٺ�x�n������۞� �u�Q�*H$���n=��v=�Ķ�'4�#-&N~��Q�ҝ��i �NN{j_��qڧEx�~�A6Ac�;{S�uƠ�:u�w� b�0��8� v�o�Eot��:�Y���#�gQ�yX��R�#���G�z�}�UGĜ��c�ʼf�C�dh��:j�?�בC��Ǹy��^7��Q����4D��7�?gcƞ&:��o��v���4�5� ��m��r����Rw7C�񯸴��f�a�>���p�+?����{� p��N���]�.d��IZ���ޛ�����(��2'+��d��+[�7�5])�Ѧ#,R.r����%�3�!|3ywiu����F�y�Z�SE����˿�W�+c�w��a��r�;j��Yo�즿���.xS�����<A�kZ�n�w���n�iv�;wp��W�_x����紕��c��8�?�����Iff���� I�=:Zz��澆2��V�*�!0j�Z���nq��=tV^;���ϔ�X�*}_�����mg�5a� ,�Ry�OO��Ps���Kv�+g�zǃt�j�ݞ�����W� 	w���G���l	��+_@���� \��\l�ѷ��:=�s��y�/�</���$[��,�͌(RX�}�W�g�e�x<i�&Cn��`�Fў�<� G�Տ~�B��H��m�!b���^kȵ�XkW�u$���5Vr�ʺ=o���/�v",o��c�+��qq�hz��F>� v#�����¾?С���.�N˹���zן|b���I᛽7Fe���11Fl"tbs�N?�-BRV>x�`�����{��j�|�'���j���ܰ�=jP��60A���r
�t�#�� �Zr�1�Z{DUBrB *5�2����>�'���N�C���jf��f�-��T���C8=�u�f�� ���i#�ǜ���R5��ɴ�G��S����?v�}@?�$�o��#��=i2U�)p2q�S<��w�{ө� ��G,��R3�E�t�ۅ
}��n;O<����xϘQ��P	ܸ*)#�G�*��F�=*�#��~����v䏺9�=kC�-f�3*Y���?.ɬ�#{��mIϯҍEt�T,��N~�:��g�5n�{�>�֝2�ʆ6�F�#�ځ�S����#�@�w�D���B�:��p���ߥ7�@�,?��@������?ʗ��׿�6��$���N��p88�z #�o J@��$����8� m�=*)�y�sW-��B�0�[��6��¹�S��)#F�@�О�5�ŋ(�)#�7u �EC��os�ց�,ghʟaMDo-������I$�.�,l�܃�?Jh��
!�$��>��$�2�OJ��݂:��� �>��g���#�j�e��� �0h�	��Tkn��^��4�t8��қ�� D@X�ЄK���{v��ȸ
O��YN��� �L��� �[�%N�n����`%HA�9�ҙ������4�6��� �8縥���Bі�d`Ƌ �\��������q���wpH�l���� ��&�kY
ʌ��0�)t���f7ȣ�kTj������8����� f�ndf���������m��P�3�.⼎A�ުx�^��N�5��o�M�x   ����px�iQ���t���b���Fݹ��A^���4�nOJ`?hl`�>8C/�ܑǨ��;.����7���af\��<��6�=�ң����� �����X#.��GpA �z�ʐ �1��Q�45��֗��r;���\<���S��C�u/��\u�$�[�m+�0 Ӷ̨&�'��["�[,:g���<��T1�6Ӹgw��/�!���m^��n��Ri�gaצ:��[��&O)��e�:{Ӡ��dk�6q�9�
�FW'9}i��h68�dԛ^V\Q�q�S�8s�@�^_^3�H�zu��)�1W�@�����:��'�S��!���Nh��zg���6�i��E"vЏ�U�渙�}�@)a���҅f�J��Q<W,<��0s����5�m��[��S�	�Va�3�:U�]V�I����y��>��������G��U�x��T^@�bm�P���4�v��l��Jі'w�Fc���1����;�@
���'���8����"����5$�~�%�tE�G�!�j&
A���	���A���dBUy;FqN��݈U,ޙ�$��*
����7�nC�=j	d�h�7=�j�:^�5�\���
��P����%�wl/�9�©!��\��mb8�T�c��h����Ҁ̼�OjQ���I�8>�x�v���cG���s�cnf,1Z�~���6���w��@�Q\�sϽ'�z�������*3�h��J6|��M5W'q�@c�j vҽE'��>����zq@
~E'?J���F!ycY�9���3�*Ε�98�z���1�[�V���;>���$?uFNH�M5��6�B*��>܂��N?|�29���Z���8�9�k���J���4�q��}�6� �U�T(ې+�� �_���p�Σu�D&(�w3`���׏�\Ay���G�J��ޚɻp�#�t:FLLI$zV	����յ��Xq���R��7�'ѻ�T�z��TK�q�Z�@�[(�W�s��Z`:q�tQ� ���ְ�!�6�f�Ԁ�h�K%��QH�Z�85���[�vh���aҲ�9�|Ԁ����3�W4���)�N$�=W�u��r�7fE�9϶:U"�	�I�V���ԞA�EWkV�K v�q�(KO��x?^Ս}!�\`�����+^Ŷ���s�k*�x�FA9��+3m��@��Z�:\���'��d� ��]�����x��Hg��͑�����+/�8��W�f[������k=U��m+�C:�VͶ�n�JӘt�_ze�L�� ڜ�{���ձ(�OZn�����=�4�U�� 55�#���.S���cJn�����D�r�Z��D�T��ixS[�J�*�s֐X��6��sZ[AW�?��I��ΰv����x�P�֦F�P������O�G�@͍"C��0,3�⳴Xwc߃޵兗��oҘ�ShU�wj�o�b�12��U�co����|��֢N�㞸�>�ou+�Ž�J���{n۷mc���^��Ǻ?�uh����9�U���ӕ�<� �:~�cs���i Fa�ƹ�*�9�OL�ڿ�w�<	�|'�-4)-n5����U$q�#޾2k����Lg̯ �7�����t���T���ocr����� �kqme�7�8�it&��w?s����<��������y&�6�Jw.�mǞ3�Z~�=���[A�H�N��i$e����x�����R�m��[f1��5��$�f���?�O�,�e�Ww֓���;(��yb�ȥ�n�����Oxk��}�Z\m��Γ^�°t��Q���+��m�C#��$��ڕ)9^��..���̠0��I�ȱڅ$Y~�qx�ƻ�zWE��~��2��rH5��V�d�0w���ٗ�A�~*c��Q�"��{RG�5W ��B��(-ۚ���ˮj�o�����⴮�d�p$���Kḵ�	�Cn�,R,��#h<�ǥL䢍!�J�����|'��Zm9ci�1)�hrǠ���\cq(�q���E~�|R��t(� et����}oQ��U�2�ToV����z��%hf1��0+�ڹ���l�A�vgȬ�Cpy$~6����:⢼R����2+����O4uf����棫&0r�<��OV�q�:W_�ȾL$����g�w���am���M����J����F[27���_.ϔr:��1	��U\�y�Ժ���@�'S��ż��~�s�Ǌ�����<�ne�-rď�}��,l�y8�������;�\��?� � Z�����z����Sܹ WC�5I�Dq֬�ڠ{U+��q�R"H��w�L����{Tv�2=GZ�� ,Y������g8��*�$�+IT,`� ���?�T΄��8�:E�FI�s�v��@<W�zcp7p���)т��ǧ(@�~��I'nJӰm�6>��ʾ[��=�S�[hJl���� �>��A��q�����銞;�f�}:�gﲼ� ܐI�)줱GQB�;�i� ^s@<e��>�$k�6��M�~��L ��@
�7}x����ï�U�T�=�1�����s�(���y�;��m���M�A9��QwD{�Z�g|�z�q6�2��rz��ʫ"sO@*��.$f$�����+o�ή����w{����=���n~я�1 ��Y^�k[�d��lOQ����"��mz��D� ��dg��ST��$`��ڶ|I�\�L�1~�i�1X�V�'�0`�]z�ڥ\Os���l���pz����^xP��T+��^+_J�;x��Ӛ��2j��؀9- *���J�M ~w|Z�"�<u�[���%���;���W"���n�I �s��u�$�O��F';Xs�r������(�ǋwr�[ʻ�<�8� Y#~�*��p���	r�E��GCɧ�)b8�9� �UiشĔ\̇l�p9����to���,���������#�Ҳ��̙��{QG(6��h��J�}v���L�.&��}�sK4�m�Sw�p1�x�D݃y�����8�yo��^?�<ӻ�s�G�T��Q��%3��������֫G*Aܿ�4���W�)� �����ެ��=54b9�
�Obj��-�=im�ɗ~}�5¾��8�RY��u:��w�Uź[���vs�`�+ھ��ŷ?l�䰍��O^�Tb���K�;�'��Mơ�[/�!��"�$�?�� �� �����]ZC�J[�T���S��O�^��{�φ�G�|5��� $�*1�pq�O�R�� ����[a�@��2�������4'R����_mu1"mG�eX�2�;�?Z��t_�+�u�~K��2�<�޴d�W�%{�e�C0���͞��?k�Q{+3��� ذ%��� ��?�I�$b�;м{�]X�ĭy8vQ���%�A���K�/ٶm+�q�e��i�p� ~\��s����|:�O��oY;}�cd��� ��REO�_����e�X�o��o'+�<q@��ſjO��'�X��!��՘������+����G�-����e�'��]w���f�0��r��-�ך�χڥ���1r1�px�j#�X�����^�����l&��WdTU�T�|����rEx��%���C�_�`[wS��p7n�?+�<���-���<3D����q�3�^]�J|X��Դ� 
�F�N��iʢ��?*ѳ8%����:��Ƨa0��������3��K�?������I��I��+�<u泾&�P�����iѤ��B�����>on��z���wFԴ_4��p�'�D���{�`o]O���?�x�e����WG
7%��~��"��}�v��!rI��3�һ/�ú����Q����l�M�*8�&����M���V%���o�zd��s�SԾ��ڛ�v^�:z��H2ʧ��W���c�5^�u��D��B��2�nF�b�ExH�m
=�x�{��-iv�q����7��rq޾��W�|%�� ��޳n��%,�=���|M��mFݗ��3��� ���z����D6�Vh��v�q����W�29��־��ۭCMx�1@�@]�<�μ��{�2�:��e��������y�˯O����#�UNSp3�+�� ��u������C FP8@?�Q��l�\���o�ׅ͞�Х���l���u����x�h�#�;^J����Z��8j����K��Ƹ�Uus�;�0ϾO5�^��W�oAl�]���jx�P>�3��0�N��^���/�����AL�d&�pW��s��;�F��i?fXż���2O�vߴt6���[h��LI�^T�$�:�Ex�g�i���Y\0�N)64��vq�F{)^��O���N�u��z��kj
Ã�k�9ݲ��e=�J���m��_�:��D���2Q�P��U�.�����"����9 ��q�ӊ���~��Nj�H�4�X�'nw`א~�zm�_���zM�Y=YX��׸������$�lֹ� H�~'��W�<����K�>*i��[�>�E���N�0}:��?h�:U���.�r�w7rF�������~��Ŷ��> >�|��`d��G�����ڊ���B��(&���1ۊwD�3�Ӿx3ᾃf5�!�Y��H$�2�#��
��-�$�+o-B�'�U��چ��h����$���x;���j����>��b�H�dV ����:�t=�n|��J�����p?Ʀ���~F=FF{T������X�e������8��BG��>�OZ\l�3��)���d��à�2O�����5X���zP��n1@����$�&��fU�f
[	8�__YxG����K�X�`���g9��_,|�o�8a����c����<o��R�����F@X��b�Fm�r� �w��-7G�X������GQ�E|�j��ھ��V�}㏂��w<ck<[�P3�S�*�F܆Os���kR��6ҩ����ᖟ��-.����P���9�'�}��p��󻰭��wO�4��r��Շ�RV����Px'O𮽤�>-�w�q�~��z<�4U���ƉWP[g��;�I�]ǎ<�x�m&�Q?j1�A������!�Z�W��0M�UbEU�9e�}��j�[���SN���.������=Nk���z'�?�������S��2�r�N6p���&�� e�v��z��Y
!��;6#^_�G|\����/��;�<?e'�1� �{��T�4=��g�=��d��l��9��+��{�W���Yn�n4=]���U0r�<�������?��������lϠ\~��U{��4�kpx��fY�f- 9��Q�iemL�>@���9g��6�yT���8�3��w5�^T�.ya�['�?�E�Z�`Ԅ�e2F�	�01�kʕ�`\q�qY�5KA�6{u|�I"Ġ�rA ��+�|?����z��4�îUX�q־��u�S��(�� ��~6���[�z?ɁX��2���qUeR�G����o��E��McL�Re�����>�ʸٓ�Rx���_UtȤ���p9�9�+�f���F���uіF?>v��@���6��-d{��	��j�Z��*�*Fȡ0z+� �	�sR��ϡ�С�yM����W������ �j���X�g� ʓ�#��ձ����Skp_ݴ��j�9X�9�z�_��z�<_m-Ǒ��N�"�$�@���n����x
���E�m��LĪ��ߩ�1������5+}9�ډҧ�NN?_ʽ7㦟oq��<'�߫��$<���O�J�sH���ymu ��ͼ�s�Z�l���tP�x`����z�h���$'��϶qR�9{�M5�*w��y<��R[�������x�)�=}S,�ճ������w�~��M*�+˕�	iPgnH#8�\��7쨷!�^X�x'���?b��jV���B��=����k��%_�������Nf]��(Ec��qz��m?��Ю�.��]Wo$u��'��U�� �?�f�o4,�Cz��a��c�O��Ҿ x���?j{k!M�F�Â>斂�E��:n���L��i�ĳ8��q��|��V�����o��0�pn�?_� ]r�ޓs���.�.�.��/�h�r��B�ס��\�WR*�Fđ�pO�T�g%�Q|9�|3�B��)s(�m2I�^n���}c�_xu�~hWW�E�8�	�k���$.}8�Y�ˎĘ!�
UBT�⑋w����8�v�E���@v��ެ�����g12�4E2M�#��W�����q�=�d��>GN������H���,wcڐ����y�o�Ni�NO8�$/֚��pޞ�1�rR��G�9�@���
��6�$���{{ue�Ǐ\��f�/-�� Zh}�{���0O|WW�� ���N�?��a��26@�+���ҵV�9�w`d��{汩'T��W��+�
���"��Fa��NB��%��9
������4Q�Ȣn�1��8��>�р+1��#Q5����G&d��Tb��y���5g'h��]5��{�lD��9��U�c�n�MR6�1���_cx[�u�P�w�u���w�a)���qK�g���n`���ɒq�*冚bLcwq_F~՟
����4^_�dؑ� {�� ?ʾv�T1�� c�+zsrFU)�=	����� 8�����P��g[�fk��}���澙�Q��5�8��c�g�j�ȺTԞ��h��=J���ۑ���x3S𞢱�F��������ԯ���.l������z
�ڧ����k��4У~�S���_�sR�9KS�t�k#�Ɏ$%Ϲ���	�פ�hT����ci��.��"l)9�=��_�_��˒x��}�]uj���2�x��P�?�-���*��r��&��Eٌ���ѭs�6�ZYE�p�+�?���C�`��]���)ヂ1\�zӔ��R�R�8�
���!GNƴ�V�c�_|�:����GQ[~��j�DQ�	X�9Q�k�r�nr�<ұ�h?�ug��)9�� �+�Կf��4��8&�s���j�?�߄m.lm�x� @A���U����H�DW w�:W��7>X��hAD�bմ{���V�����֋{)om�p{��_e�~��a��ז���a�Tr2{�����F�#�yȯS��ߩ��1��?���ƞ��b}�3U�]�Vmk�)�z������lc�{e��c����^���d�b�U%Fq^,q�=����������[�[8�t�䵊96���n�� ܛ_�1�IU����O���x�/\�j�x7(����c������ǖ��c������q��<���k��>�iՑ�����
�c��Y��\�P	�aQ6Έ�(�/���}���W)	W�6�����i�G;D���k�W�F����	 �D�ɴ�2+�/��TQ�Muk�G.6��9'�3�d|{����׉ Ve�:W��?������`-�g�һ/��
���A�` �H���"�t6ij�s�W>!��,֜#����������@�'� �\���Zޠr�����9c�u�Uabq�_x{X�K�y���V�z��l̪�E����ŧ�����E�
/�a
��Fp+��Ϭ2��?fx�Yd��S���B��9ju~	��m�A�bPz�?�߳��k�X���_Ҿ��U嶉4���������V��-�eF��q_:�u��c����Ϥ�0�m��Z48
đ�W�|5�y&�� �	�}_����u'h�]���WW��pi$:@����z2�N�}Ӌ����y����o6����}x��/���6H�Z��8���7ȷG��00�r?�|��]Y�ŧ#A���B������aeS��&�cf��J�j0U��[�xgPxRk���h`q�{���X�Y�督��e���}���\.�+��2�J�+C����WM"KTbV���rD��6�/-�����|Y�w�־CR�;Q=�|�6G��G��7�n��'ݎOQ��x^�'�m�&�q_��;�ޕ�k����J�O�6=f�I���b��z�^Y.VEHS��g���t�5�[�wz��_��i/$P�`��@$W�[|7O��	Ƞuݟ�WX����l�Yvc�k����w�Z�<6��V)o��#����]�3��^��]j�]x��(0V2=pO���Xn�O�Ҿ�ۦ��<z������Ȯ��I
O���<��>�m�h��s�E|�n�n#e<�N:����x�x�V��G�:�ܶ5�$�>���� �x��;>Ύ��U��F}����j���$�kv�v�k��>9�t�S妷��f�~���.��<b�[��-�@���6i'f�?'t�7ך�FBT?�����[���2���<WҐ|ђ�eX0����h#�-�*�8�*�B��1g�x��}���dDG��~ Y�x�[l �7~����χ�'��.���������R�}/���������"���HO�a�q�}ӛ[�u�rǥM���g=1�+O�fkid1�$�\��ڽ��-��GY���fu��8<t��1_iA:�|�s���߂�/|x������S�$��|��!�#��O�H&_8�
��J���^���Y�"��j�m�7J��.���T��k1� L��~5ZiY	N�f)��;����[o�3�5nW, �
�
�0jԐ�@q@0�epz�5'��\ԻS�� ��<���+�=1�!�X�d�Q��<u�fo� `�a����$�b.:zVF�$���t��$x\����l����t�J��3[�}̷4�����H#I�;|�w��č��������1�=rC����1>���ř� ��Lt�Z͙1׎j�kZz�=sP6�k0]�/��i
�Kb��w�cw����a;\$��j�jV�6��{�"���@�ӓ@�	nc^{�!ߍ5��l�p?I�����ހ�����T���T+�����jռ���d��@�)hY  ���?�(E��98'��G#�����j���\�4����ԃ��H��V.���q&Ч���w̫c>H�6�sڢ�.��vH�aF���/x­�\O�昐�(���#�ᶎ�	��H��r�|V��{q�}�3M�03�s��=�W%?�kV����K|�l}?_J��r~.֯��T�܌x�X:�����y�)�b"@Ozn��Ŭ^17��;�����k�zO�pY�ӟNk�1KTc+�c�x�Ě���G�[h���k.��������Z�º&��hU ���*�Y,L��z�Uila����*;��� y��������`��a�]����½O������IY�G��NFIO�+����þ0���,��y`z����%O�c䙼#p،�F:`���y�6瓟�_Gj�U��"a$ �>�ϩ��T��'8���d�#��[6�*���@��Ҵ"�/-�P����`�׊�W�^����$7Aa���ױ��ᕟ��;Ik���0b������9�e%dG+L�"��]�L����ARG��Ae�u�	�˓�N0~�W������k��l���H'���ו~�^ _���tu����qj�)������n���*Z3k?/-�0Ň
���K�5M:ۻ���3���+Ǔj����������;�%�Љ��>a��\d�ȏ��F}Į88��������?�\��8�K�$K�ė2.7g8$���F�v�x�&�Z��t7Y̓ U�FO^+ꯂ4�x5�ˢ��}��|�1�)P@��W������;�s��<[���>��&K�ĳ1��{��:���⫉mV_���;�r���e�l
۸����=��W�88��>�}�|z�¿�t]��U*��yP�,>�i���o�xP�����"Y0N�� ��Au*Ŋ��jE�' �޾�6��п����O��z5�0[ͅFc�{+��{7��E�� �7Y�{i\��w�	=F1��Q�+.�1����jo:�0��11��wި�Y���Q�K���v�u��yQ1�p'��k�ί��[�s� �ܫ?
����  �r=qI��2��)����~!~�W؍7@O(���lg����n&�R����O:�F�����M��n��7zw�#�~��=)�	�%��j����I�F.k�>&~ӷRI���ͼ6�|¹
r �1_<ya�����5�&`��Kd�����Ϡ>8�h�� �M�5ݤ��v��>�����y�W��>����=B!�u'�<}}+�!_���n=��uź�gU8?)9�t�&�d�{�7��q����������' ��_FK��@�=�N7�G4��8�i���Tu�2o9��T �%�:� �_L�+�V��o� cꄠT�C7=+�%m��!�})�t��*s�O�T��c�|L�����3K��H���#�u�s���~��	'!����}OʼQ�i�R��y��קx[�z���LCq���j؅O�6�I�Dc���� ~&n�`��U��c��9�@Im�P��mnr��020O�P�|��{J�� � ��!䋟�� ���4q�۲:%��Wg��q��[����m��O��q��=��߈�._����(�5�z�δ5�	��Ʌ$��^@f�Ƴ@߷��}k�K�\���1F�p}8�q���+� �#4�]�͐��8��9m%P*����IY���'5JAk�[�kX�_����i?�I!���w'q8�秭y���X� �uɭ ����$1'�� >��{tΡ������o)�~`C3T�rTluן�o�W�"�ܑI*���|��>��z����|i����8��Lx$�1����u��V<��G6�������v~(�t{I��e�c��>ٮg�g�+9|.��Ln$h�v��l�W�æ3FQX��x��a�$�~~��?7_z�},J����TbS���ni 1�?Q]x����
���[� ��֠��,[%A�9����i bk��њ5`�2�v�z��/��?�(�v���җ���9�準�V,[Мq�T�<J�t$s�x�EЌ����g^���bH�c+����4oxr}VH��3��������G�UM�q�je�F�æ���E+�1�?>+E.���Y�f��Tg�zW���H�� u�һy4Hd�-���EA6����9�<u�{�eb8�X�>��G���sڹ�-/m�!��W[!���?*ټ���B�=l�c�:���,���\���%toN���~|j��ԏV�V{s�0N�:u�����P��-&�V�������Eokb��j�^8�{�Y���_gIv+��^ML�Q�zP�E�����t�G���z6��0��� ��1�<� W�𹅙��l�rrG5�ċ[��-�E|�G;pߦ�|�!��tn '�<.!�#���}��>�Ҿ;E������n���0�G�k?�{����wksc};Im��rO�^���!�ߞ���#[�<�u�뜭\�.x�O��5snēlh���v�S��W�"ı.0�Zv��}in2K;��n�}�CdpA�_b�O�ƅ��Z���P��UFW�����RE��G���0B���o4ԹD�ϩ>;�X𽧀����"���n��\��x���A����w�-�ڇ )��W�� g���� /�9`e'$��:R�bQH�����|-���G��;�d������#s�5��RQj��&p�?.�|����#��<Ƕ>>A�N�S�8�}����K[�d�h�r���g�x�_������ŗ�ĩ�n$����v�a�w�I^�l����2��
N��ƕ�^`#q���˵�B	�ڝ�h�/_��
Z9#4�ϧ|�~�Ğ��:��lU6<��`�Ezd<)�����G�/$���R:��5�h��R2g�i����d��G���|ڑ�}#������C$���G�4��9Q���π�/<�\�܇�ӱ��y$���&�T@cn%q�R���m��7�ڗ� 5��k�e^�8�]�\�O_S�׫i�8�*^A�]��%�rI��zW�^Z��E0ڝ�=I�O�U͠�O_��>7M�K[��Ͷ��/�4�2I��}�Z�xAU�㏽M�&0����OʽEM�Jü��ɫ6�.ୃ�$TV�I6�Q�s��QۜІZ��?�� c?�ޟop���.0����^g�ېĒ�U$��j�0M2FI���8>�9�8b�p�sۚ�ݸ��Z q8���
$n8<�=��Us�T�cXW;w>:� i�/�O�Ia�3�ֽ�fI�4o�E	-�#�����I����}��n�t�W����z��ZQITbe̚���q��Z���Q���=+�|+�1�_i�q"l;s��[T�Y���w4q�9s�W%�k�v_|<��y��DS�JǙ�kk��xW�����J�'ᯈ�l�x�eU�8$w��<Q������jGl�H�W*�x קhz��V����	�%th�>���#�1� ���u��K�nw���+���ռv��s!=��_L~��u�2B����\�_���Gg��p����Z��=%��<�\�L�giåX����W�|F�C0���^�w>'��5����"���|�=/�UQ�y9'�� &� �S}���+�C��Rh���l��g-��s�_�W,��wL�����=+h+lgRM�Y�S��2{W�� �v��E^����f�EG�s�_M�W��C�?*jEKV:M�{ 񆳣��9�vH�1�{���A��	�����q^k��Æi]�=��S�
��V1-	l�k�&�GS��>���G��^XT�ޕ���c��$Q�x�k�z��.F9<pk鯅>,���FDvZ���R��x��>�hZ\�c� $1ҿ&?i�Y,�*��� +���?���qul<3y�20(q�k�������Y�2���9/�?J��ry�����L`��c��^���mC�R���8'&�H�4���VA��	q�$S�����c*zH���ό��<27��b�� �S|=���Yu�b����n��q^V���@�2l!�z��_ʸ� ��NY�Y�_ČכN�����_h�v�'�'�X����^��_ثp�����/�?K$�ZB�ɯ��;�e��8>�9��[3_tt>(�Yڙ!v�x�^��oU���9'i�z��u��?�=q^�f�M7N�����W�^��&��5������ ��Sp7=�����Y�!�A8�kx���F�ǔ7��̙�����ʾ����"���@�Cv,��N��zs_`}�]h{n8��|a���T���܎k�&�2��`3m!z~��(�M����k�]H� g^�֯�Z�a�k�o|Q�O��7;��ҟ<h�%a")(��{sR���(��;%�&X��zW��Z��o�Yy[�O�_Y|9�>���T-����e|z�֛��tG,wn^q���mY�~~��0{��D�,�1����#�8�}}U��"�Rr�d��[�m�b��ʮ�H�m�%H~d�=�_B���b���������	�޵�7�� ]N6�)����F�w�>���wz|c�g`{4�;⤒I�h��f���_�Eo��%H���WK�v�g�	#h�4�*�Z���dοi.���:����P��y��_V��_t�f�[��|��5�?������Q6<�/pp@��U���|]s��y��nldp���8�����[ӥg9�+u=G�?|=�����\l"9����nxv��:���u�R�Py�c�����Q�3ÿق��ㄡ}�a�ЏZ�y��<h>!|D�u8P����D���1��׃���WV3�)4�>7_���#��
��	*={��H������b��H��ƺmuc��g�� <J4}�gh�����ƓP���[ �͞ ׼��~#��+Ӯ䅬|ȎI^H�3����Tg�^	���t����g�}柪�^Y��H��Ɂ�h�~E|=�Z{$��c���_a|1���x=�[��7�\�zS�9ZÔ\�������j�[�G��I$\ �{�k�r��-/���*��J�|�L�<y��`�����5�ω|3>���E-�,Mi�Wf}Ϳ�f���/�,�_����B��J�ڊ��U��T+dp��?��+�Cq�ں`ӎ�5"��߲��g�z�k��y�խݗ=�k�:Q��V 2+�|'�%��C' �f�l8+j}5��~��I���=NG���qܾZK��+��|`�÷��ܰ�N3�}��u? ~"�k�e���x^s�\�&�s3��9�I���]>�4r��I���}+w�}�����%%E�KI�u�SV����������)Z�s���h�/�TΊf�2ˎ�{���5��A�{X��nARB� ��~����*i���5�3�ٞ���s��oM����i�FF\�]՜�`�kb�h�-
d ��5�ٳ4��gڶe�1��~Q��+���Q�2����c�z���.|�B�9kr˝�����VI��������z�N�J�.�FV?`>�R��	�1Q�'�YH|��9��˯�O����t79�]�w6r3����y�]B=KI��A�5�����-����0�8��8�;�����dz����ǭM$�n��ڠ���i$c�� |�s�{��o�����ަ�ܹ~99��ș�p�{Շ� V0��rqҫ�;n�����ӷ�i\뛢���W��g���tF�B����N�W�������⇂d�rE?u>���[ㆧa�c����������&%pO'�+�oeyu	7oU9�
κ���1�/~V���mH��,O�Z,�b��������N�^�'�9ۙ$�q#��V����ߞ�z���38�iMc��䷽Z����a�f�WA'�vy����e��S����f$���7g=��]����R2>���?��Mt�r�By�޻[��L�ٱw^�楨I��m� k)xI7g��o�Xgj�=s�lj_�-�e��<co?�5���;�#�Ǡۓ����
�:��Ы�@��3��+���쳔�g�}+����/tK���;~ꃟֹ��{�X���麹$��6M4}��C�D�ѳ�c�Z��Bt�Ն��w��� �_1|=��ү�B}8���7z5-9X��G�J���K�;�X���|�.1���<��u�F(�
,�&gi	Ǡ ~�k���o�iL�۞���jv03�[H�If�i�c3�j^*�|e}5�Hm�mQ�;s[��u�G�i}��E���#�Ͻ}̿�?uZ�f\�*	�o�����
���Z���%x�A�]��){�ԇS��m�jxN���rһ����*ms�d��F�GxP� $�f�|���%��"��ߜc$�Q�W}�x���z�EIxr�N*�w'��_��|3�7�^%Ԥ�;[7`��L��Q�_8����ωn���KvPX��#856��?[��O.\Yn�J�q�#�j���;�p�;�rN�Ã߮3[9s�Fe�lfi�<��ڶ����
Ie�9��~�I�#��P��>lЃ�/q��F�ws��|}��K{�d�9��Z��/�Gº�����[���+E���#��k�ˏ���_.DW�z�4o���� UEOa�Z7qs\��w�ڮ�とZ�1�w����~��7����~,|T���潶���rz�=1�ƾ��O�<?���֤DQɩO������5�����5֪�f9f.����5�SXǩ��o�2Y�@���
������}�~h����YԬԴK<��:�MG���\J��8 z�&>-�� �A~�u����jS�`~S�=�5��Ԯ'�?y!`z�k�2�Ƕ�?Z�Ǟ��W5#}�$`���Tj���G��"3�`#-��T!�����zjhݸ��=d1�J����cgiƀ�x�߽(��9�jn� S�]ŀ%q D@��� �G���q������B�9���Re�L�����F}��;��;s�68�RB�簧�0Ux����,���� 
O��sޟ��;����}��+.2� 0��>��$?*�}}jF�-�g��JO����g�^h��l�+��z�X��:�Q�<v���wh��A��E A�� �A���ݻ��� v��M=�l��d�f��afW\�S1��>�{����u�~�,�~��ةa�'¾px� )ګ�p7 3�+�[Ųiz}�&���9�?ʼ�M�}���1��	����o�Ioec@���5����]��3�f�����*X�퇬��\�|�q=7��*�Ǉu8c�S wX�Mn��S�~U�O���6�k3=�|�ߚ�kVo�pEe�� �����M�ąN܂�ڽt��滽K�gx���4����}�H�7��e��_��W�ظ*0��Ӱ��4��H�#=s�T�`�T�==+��R����d���8=���YH~�8�:��ڤ�=j2�����={W>5k� �:i?�.I�$�q��`:���oC�y���g��1��R�ܣ+Ӟ���o�\	-��� ;��ߌ����gMu�H�n��Au��K0�	����ܴ�0���:�E���u���xWr��g���?G�X�}1\�����X�ZjZ���������D)�����+]E<��?9�'�ɂ�@T���nX�2GO��~=Z0����D���n��9�y*[,��C֘2�����ߎ��+x������r�F~�8<s�H����y�H,tW$��mU�j%�$�hF+��X�B�t�7 t����ª�>��X�I��axꉗT�5PY��:�t���,�7?3s��X6�|l�0'>�����UYbZ�熌��Wq;jMq�X��#�돡�x}�f=M����^�g�� m��l���;W>������f�c�9=A��=IYժ�G��
�`1�c���<���{�.O��m�3�OJo� v�����k��<�3�8��$� �����A�hp��m������8�#'�@̶S��޴��Q�p@�l��֡���Ӱ���To��~��C|�:���*�_���Z�aEV8� ����U��{E�c�� �OJUa#`�ⵚ���x�*K[Xc�����a�Us�l��#+��}��1�s�b��V@R���dUhbw�!�浚8�0=�x�F�
�rwrh'S?T҅��M��p�K��mudƼ�5�ƙ!�jױ�|pib�cحՏҀ�����vd�
X�'�U�9�zW���i�ǹ�9�Au�i��mU뎔�"Ү&'
ߗҖM.�H��]d~#���.j���C<*� _?7���=�x��Oo2��m�Z֚��dg۝�����92�{�ZV����K���܎�����ԭ���;f���wU�oӁ[zo��4�6�^�7Bh~B9��������\pƠ� ��7�w'����jM[���[�^rY�ON)���s��1��Z��Yq�t��o�ޕ^�O����,C�dp>^�55�nm�Ӎ���y�UU�O$`g��M���C��|)��յ�D��� �A|to�����h�"0�>�J�'���v�E=�m����t?5_i-�,V�>�Iǥ=�5s�m[����5�g3�h=��������!�l�F��la��b�f�%��u�7��`kc$�"1�sY8��M�Y����Ȅ��� �� �+�����W�pOOj�Y&���C��g<��{���Z�M��'ڕ�Gm��a��[����e�V�m|�uU�ܜ_3���o�"��!�k�~�.�G) f�z�w�Y�[ݱ������M�����>�5�����dѦ�"{sT<S�$v2�lT2R��������K�:)�!C�+�����_K���u;���Ebvt%��������i	R�tEhD�M�S����n�k'<`b�j�fk�99 ��_��!�:zg56*���Z]K^a,��~�j��O.�P�S���+�|u��z8�$�	�>��r�Z���LZ��7����]�t�wV>Z8�W�|?�f8<���~��{��W���c���l�՗:���\w=� R�'�����Ӂ�j�u���Z�����C,�\r���\�u�]?òI3�F��wl����q��|q�r�Z[���0 � :֞�%{��xt��&��ȭ3�	2������b�����W�.7�(_��c�u�c�}Y���MA����Bc��esǯZ��_��4'���C�Jͣ�三IH��rlΓS���Rբ��"I����?ʾ���7ZM��ۿ��~=H��� ���+�]B���i��S��־��?�=���z_�Z��F'�1�ؕ���g� ך�RI�����7cV�w_�g�!�@h����ڸ ���>h3������I���sߴ����WE�Q#����N:�Z��N�	rJ��o��jAGR>c��<⳦��[�q���#��5}�����Z�����u���w��)�>6t�۩F �c�dW�x�Y��J8^���?�I�w�cy6�u� �^��O��xbt�w9ղz�ExX�Rg���4.x^���q�����ӿZ���[�%���e�F�O�:�ƾ�e���7��猎ٯ��x?Q���!<���S���9�Bͣ�]sZ���(�$V�89_�t�2M�hq�b�OS��&�Y�-J��}¾�<�t�dլ_K��z*�IǵTޗ1KT��� i��$֦����3_�رV#ߓ_p�՞$�='TR��@�~������b.-Y�?�q�<f�'4�*�l��m�=��95��W�S��;H!{�?�u|۫[�� z�<��OٿVm/�1)�,��+�Z�zb���a��ㅎ�Hԭ�_3���z�g�\Z��Ã������=s�7�x�V�!�\�=#v�t�+�%<�$ϵ�#�<WЖ� �񂥼[D,��޾V�O�]c\�5�;>@�b���{�>x����\�A ������*QH�f�b�t�U�+���#��ϟ�A]�i�Ry� ry#��E5���Η2H��9���'����<E{�����~�)�i"ct�|�џss�c>�*1#�º�=	犳���w�z��v��|&|Eb	A�^��xZ�E��@8 �c�s_�a��eUd���+�ZjZW�nܹ;G^+��I�p��߂����fy�3&r}k��h�A�"�~�_��c�UY�+c�}��w��z��R���W,➦��s��k�=��$�q���[��%��W�YCl$0=�+�Լ��,W`^߅|���˦������G�zqYT�k�-��|�Kj���c�۶����W�����H'��b���O�/8߼�$��g#�u�����J�N
�5Ys��|	��Eh"s�����L���,���|���uH ݀�����|���ha�Fy�yX�Ϟ|o��}�L�un�8�U���Huh�e�s�g��~����rúP:�|?ռ�5�07��g���Ma5doMǚ��^�5+;6�ӥ�or�H�W��[�&�K��+��z_쥥������ƿhTE��NO�ү~�zo�t�9��w/���yǩ��.�Gs��r���=�shG�K��
����u�� js�Ύ����A���'��]-��4�N�3�鎧5�ψ/�Z׮/vL��'޷�NU39��0�	���2��I�]6�,6*7|��+ߚ�->�B�զ#h�'+��9�`�#�cnG�nY�$��`��Q� �u�c�����Ɩ��ͤ떗�H�d.Ї�s���_�� ����I�7-�(����q!en�pFp:���b�6��\ρ����sXT���~�0����sL� �}i�}���R���#b\EgbG�N�,o�pEG��� ��㊐>u���6��"�]n�eݽsۚj�P�p�Kr6�$׈zD|d��ӱ�$q�yQ��L���ǟ3�Yj�j��<��}iג@1��T��� �@x��S�����S�=�9�T*� � �/!�r�:�Q$R�ݪ~Y�q�K��N2G��K2�3�>���w��}E=���G&c_CN�z!h��
2=*f��\n��v��>�Q��:�ސ�yd@�}*��� "���Js���֞�y#��1ϖ��X����[x���>��G ��O����B)c�+VB������,耞��C¾-6(�I�z���l�+2���\��� 
�lf-#dm���f~gC}p�^L���H[�&�56io���6�c���\i��q�C��U7���k|���gֳc;}<;["*���^G�Ki�xn��wo�L|�zW�ir`��]�kξ/^C&��,�A#�~����"j|:��5�:�֏�hAݳ<����[�ߴ��m"4+)@s��\��4�/*��F���S�"�[H�d�q�޽��jy��3޵�ڻ^�t[k�E�Ȯ�3� �E]���u�
#�@�nb}1�W��� riWlq� �^*}��i�Ϣ���.���KTy�e>�{��k��� j˛�5�6����>y����~f� x������8\`�95j�E��Po��r(}�X�	�?ʯi��e�]��jv�R�ʼbE��z�i�ۖ����A���bJ�?H|3��	�|���j��	��ٜyJ�Hx���_(G�z�ke�2�ۻW�M%y!UA8��?Zʒ�-Po籨��SOh�c��*^\"�̸���/^x����H��T���qy�z�c�MB��T��Ha޴PD93I4� �2ps���U�4�?h۱� ���ss�+`F�����+glz! �Г�����,$!x���X�Y��p|����廐���W'#��ry��\H��>O^}�5"6� ��T(��ڳ���G������ۮ �lʣg��Uh�g���p�F3��,		 c�EA%��C�d�9�c<V������zr��@�RrQܸ��c:8"W��z{,E|��^�y�;/���`/_zH�I�=���k>ti�P[X�M��9����h��d�B�[o��_�0ᛢ 2h� �]�.�X �}����/c#=��� .;c�ME�X�s���U�;.ޥ}�:�$���s���S��~�E96��?N���.7n�H9�1�������i��tn;8n@�x��{D?c#!'H�wۿ?�D�d`�w�q�9�+}�82]Ww}�;z{V+���6�Ď��n*�+��#�h[��܆i����J{+u$}7S>�)��=hbkiw�.w0�1�r0j�]D�w�߿��>���z�P�4��|Ͻ��r:�q�.��o�PY�m�3��]S⥢��ov�xϜU[�0���n,ǟ~ơ��dzM��כiE�����-u�fy6�q��F~�+/v�$�I�=c��֝��B�)f��z���Y�H�#�Ms�FA��Jk��Iq�u�$�����S0s��S
��=8�����HW	��?Z��V^@ݜ棏�'��4�6T����Ȉ	�{)�/�01О�_xP�=�?Εq�קZ ���Q�O���c��r�'�v�֫"�A9��4��
�$d��h����ӡ��S�a{u��JEs�u#� �Ma��On;��wP9�H�}⧞���f��BAB8'��O�S��Uʠ'�R�e���F摂g��z����9 ��hl23��z���?0;����3F<��=i0�H��x�@�W�ޙ8���^����P��q�����NǴ�� C�'zt�����|"@�>��3��Ǘ$g�ϥH�<�ypz�P��_���X�v���|ц��1�'�+��c�p(��3�������~166>KA89�/�&�Vl>}�W
O�0O ��$��)�v����&�l|U#2����NE1�Dꌬ��C����X珥;;Uw7�Џn�
ķN�;1a��OZt*]XFN~j��#iʑ���*He��'�)�=>FnW+���$�������\cn
���0�y�ִ��@�=9>��d��t�+����˥1���['py�]�[vH ���,�)[<`s�_�OΗ3�G<-ߜ�~S�M��߱���	�=؋hC����Ơ/�I����sW2;ҫ��<��U6�X��s��Ҽ��v�}k>e9�^sZ�s��m��A4��*ۏ?�7`s�/����'�F�,���0y�\��m���MTY�c�/��=O�E���e��>��V.�1�x�ZFo�=9���9�_j[]���׌q�ޠ�F�X��q��ޣf#�0=)�&�zSu��8��d`�s��u|���әLm���C@hhi�Oj�0OM�鉚b��^J������u� @�h�/�X濆B��a�0��Q)�ַ��%V\���f)U�c��׊��M���)l"
$�nv�u����S�@\��� צ�t;��RW����/t���A�(k�UT`��t�"HHU��4�#R��T�*�Î;��f�$pc�V5De�`:v��QG��u�H��P���s�]���Q�"�Y�ϯO�5���>�_hH�;�v����e}j�y�!Ws_S|\��4��8�YX�D�NIc��4�f2��<z��]���Īwzb��~�:u���c$)#?�����/�2K�*!9��/��R���+i��E�5����.s���|3x�D��8,�+O��ڢ�|�lgָ+���&��>����Umit��9~eݞMc#t�>��^���H��k״V��~W zW�^���j#v(Tm���Z��n�˹�A����4����-:���z�^7�#ⅽ���T�$���ǭCYԈK�D��\�<a:$�wW$�*����kv'-;����wXev���Er�q6=��V~�4���NN��֠��}q�
�S=�5���'<
�x��MB���Z�pMx��ڿ)/������œ��K�֥Ŵ~�h>&��N��W���R��ŅȒuU��u|��� �������v�?�h�H�'P&�f�v:��^�y���Y 潯C�+%V_��^��&�o�����k��G�U��vR4,�c�Z�Qm�s�?h_���������b+�B�V�y}/�$�����WG�g�^��3Tv��Z��(<����8�2x��J�uf2}��M��A��3YZl��RG�U�Ͻ1dc��}8���M'mt�s�w�c��%��y�+�t���e�q6�0}���{�Ҡ���O�'��v�\��i�6�����
�ة�X���������P���_¼O�����[���1��,7�¹�'�������wo(*�}��\R:wG�ZF�i�.餎�v8���m��KF�÷���V���&t9
9#���^�K����H�Cd�DmTR:��T���u��;���`�3UNv�2�Vڐi�
��f�<����i�樒�
nųP�����T䷑���7��z�G�w-h����[���������$�vЇ9�b�8��d�5����R��$����?�X�5��B�����|=�;5E�Qv� p+�xV���\s_�������5��p1�pk�to�������z�R�[^�S�?­�i0��H�~f��Nk��:|j���=��*,��O�l���#������;��x�>2k*�X-��),{�8ί���i��J� ~ I�-y��̶Y72��q�e��P�[�a�Ɔ�X�vl�#}��Sl����q�kӧӍ��9Jn�~��K�����;�W�x3PM���vЄf�͡}Ǎ���5b+���1�S���t&)�}��� �ֺ���J���Z�|=cc��;lec�{��G��RE1�i"�C��5]&5A��� �Y�������^��t}.?!ڌÕϮ2?�};uq���N�1�gi
�$��
�V��xN�n"ܓ�̜���Z���� �ǎ4��%�|�9�@o�&� 
�rq�Qn�;M������K�il%X�"�p��c�T>)�]��3;4�hc���[~*��������? �>O�z��7�1�'4��q���
�\�c���*�3��X��cr��t:֟, 3���lb��Ф�T�xY9�q5fv�	�i��������?>)��lv�2�۴d�W�V�e��d:�ӼM�h2	-�a�ޓ�f������M�5��2�?J�?឵��^��y�Tc��ˏ�֚���V9U�����/� l��d%K��:� J�)��~d֧�/�ߋZLzl�.�fU������G|]K�n��ɐ�(<��_ڃT���ـ<rkŵ-B�[���FnN<VT�������1�J:z��n_�I'q�X�K�Zk�|��LS�
��8�Q��8� g�zz�pw���TWVF�8� �O�_�(4;{t�� k����`�jh�h�ђ�CUk���?�g�� ��cY�Pǳ6k����w���0��N3_�~���a��L�y8�z���;Ķ���p� ���R2���q�Ͼ�?���9��m�` �)=@�^y�g��ǉn�� UԚ��\*�­|�y�Oėć��ճ\�����5�|�u���l���KCS������>�;K/�^]kl#ROV��k����I�ǹ���O�73m�!��ӧIAr���g�[��X������"�~U�	�����{0Sojg�� ����<����q��PmP=x�R�/�I�xD;���N���~�][�>g�⠸�Ԗ7\��8d~�� h��pD�*��V�������jд2�[v���}~��G�w��CXB�p1�j��vq�!s#��u���*�ڔ��ێ�I�s��C���Y���6�jn��r)v8RZ��h��o��5�UOC��@R0@��r�$�8��r��*@���~1�~���ϵz/�?���CBm�`��v��<�c��8#�o���$����ald� ��\�)��h�ɟd>+�=�J��iA"��C��m�Yd�A�2�i-���?���8���d_�T,�`� ���<���k\30'�EJ����֥�5U�Ro�;�S&S�qޥ\� {�|v���� ��Nq���M�O3��|�� `*2�r��v)4��t9�d]��:Uֳ����t�����3Q��z�b�@���?Z�a���֦kEh�ڐ��c�$pk2T��$g���-���Ӭ�n䁸��)?Đ�� �Ԅ*���N��r�_)�� ����~2��nW��z��!���00Oj�6Cq>�g�*9�n*.��}��:sZw���#���}#ú���IQ���q�B:�Z����y�2���nմ�퐣`z�� �������?!*��j�ψ����ڴpI.ｰ�F+J+������p��1Fŗ� ���̣������^�5;�K0���"��Fָ����b��.��J��%ec̔d��������V݀?T�*#��<t#�V��h���$���\D���~��wv mє������T��£ך�i�FG^�>�ֳ��#��8�TA��3�#��aR�)_�>�֢�6)$u�����Y/�ݎ�56�c��n�F��|�}O� Z��B�n��6��&㡮�Xѣ��cixQ5�@[�q��^Z�W���ߥ#M�f���H�=I�j1rV>>aԶy�#bd(7cw�� ·>�hE�,�d�	ǿo�����j���'9�Ա�]�s��Ȯ�x�r}�I���z�
Y��ھ�j>FA�Hn��}�H�G� Җ��4m*2	��@���#p��ֽ�>�Y�ٻ ~�sg���FI� �פxU�M;�݀�;{��Ⱚwa��fa�&�d��5��¨��h;FX�rS����
���@��!�b;dc qۥ5Tm�����R�|���-��FB����U� �r~\��ڒI7��m�s�U_ݜ��H���1��L�#�)��Rn���q�Q�3��c��KT*��66���~0k���y8�Ƹ�E�����tS���2l�sߑ�M��c��;Q�lU���J�;�#���8�`;q�Ǝw�T� ��:g�hV����ڧ�ǭ0 ���� �S��9�:�g��J@�{px�)Ŷ��*���7%��N�G�t�L	Bʣ[5��9����3��(m�d�H$ O�,g����w?Lұ*H��S!�?_��4�܅ �g��������q�\�H���I�Q�#��>96@�ё��+K�)��i���8�?#n׭65 ��sBv�ۯJ z���=K���5ݴpT�~��_��O4 �����O\rCc=*���^q�qR��2۳���� ���v۞�����z�M�6�8$�h��dgӀy�G�Le���K��j6���ӑ��nԛ���M�}i�D����N%o�C8�=j1�"��<
Y��#��26���P��>:)�JL���3���U��t�g�73`����(�:����I��� ����RHS�3� ��v�� .ѷ����f���4m�	���i��PFFv��O8��k�#�s���C���pA#1��J `�����◸P�
���x���Q�7��4��L���Gs��q�F��d�}_uϘxU�:��#�������dv@� x2�؎��\��^Q���=rF��Ý��z�ʢ0��#���Ucg t
6����HV�~���ը��ǌg��l�X����Ҁ�s2�+d��5Be���G�Z�Z��X��g�6X�����yħ�`�@=�9u��.F��΢�A6�x�W >�3J�O$~4��$��0q�\�P�$� �ɦ���Z���@&��֤H����ԡHf&>y�*�w�[�?�#L�9-�ֆ�Yr��F�>��@�y�T�������e��;F8�>�����%J��޽�_u���J�8��8�$꨼�j���;����1�����1��b�^�//.�󦜖fc�$��YQ)�d^�1W�m6�N��␭�sT��g��4��>�-p�������l��|��/�9C�ۑ��tz��m�f���vL�N��>x�\�� U7Rm�D��z~�l˵��٪C�v�.��q�����1Y�$���x��7��[�!	�=�%t˫��ag�*4�.敂B�s�����+&�X��,p����k5�������型?�^9o_��V\�m�hϯ�I�27k_]Ó��t�^��{��8���eɧ���:᱕l�zʈ��tPzֆ��Ԯ�Ò�=Mgn��?�[UU�05V�T��E�-���`��2g<u��T��y�M����k��G��+�̣q'��g�/��l��-"Sr�q��ɤ8������/��]����4��z��V�X����>�!��w���_Rxg��p&m�. �Y�Εh��� �u��b#�嫱��7�?�1�"�J��XAǔ�������/�V��s�̿�f�� �A��G�,�p�H��~����U�1��R��,s��q���5Q��1��:܈C\ˏzs~�7�*�]��_�+�5x�P~�� ����_ʧ�=����sxA�TR~ɷ`���LW�w�":��_ʣo���!U���y�Q~�w{����U��-�m��dt�k�i���ac_ʦ�Q������<���?e;���a�qZ���C�U?�~�� �+bDk�R�؜�-O�G#i���,߲���0L�Ƨ�����̷��W��fǴj?
_�F�ƣ���������Rڀ< �{~�g����=~��
-*�~ϝʿ�/f������)H�x>�(��G����� ��5'�M� �n�u�*^̞v~{��'��@��� ���h��C�ӭ~������K��e��J�P�g�̟�2�,{⦷��m�s�� �=�C�T��U�F�����,?��m�7������U��WݣI��Q��j���C���=ewdD1�E?�N#��Wݿ�6��Rc��A�R�b���T����q�c��&��F?*��t{L��*_�N�Z�T��{F|4���A���Ҭ��(ڶ�����k���mG��S��m� �����>?����� cң����+�A�|Wܿ�v۾��T>�h�F�G&����_~���س��<W?��຾���1 ��_�z����Y4?�x�<��~ז���s�M�^��tϖ>3|���$�8S��WΚ
�e��1�(1�
���ώ�WI��DY�}��� �������$��Mj���|��GK��5	��8����,d�[��������=�j�S�o_�ެit˷�I"r8�ޯ����'��֛>��fVRǞ��[7�;R=�ǵ}9�A|�F�7���>��K�/���!Y��y��X��\������a�#��Y:����1�6	�s���0�	�[6H��x�p���K���d)<h�}ɍX��=#M�՟ˍI?C]N��W�`~� �]��]?O��2��B�����>Юt�&#|/P9��S	������R�������-��K����	�}��r���.�(w�[Q�� �|Q�R�'ؗ�[�}jem��]��.!x�W;�8��ҷ�m,v��zס�x�O�ñ0P'�/#�+ȟU�D�c����rߑ�i���ǿnZ��<%�"����d��c�=�]g�/V	�n�Ɔ\{�����A��s����k��-�]6fU*����ӥx��>)ǡ�@�ʼVW�ߎ��k�K2���w�I;��Oٯ�:^��^�1ĊQ���z�~�8�g���G+m���_���o4�"X���B<�s�3�s�W׶� �k�&[�eU$F�0x�XTNW4���ɏڣ὿ýj� @�� �¼gC�*�*6�c�5�O�� ok�RG��)����� �&-�c�χRU�8��?Z)�Aܹ5&�n�ጺ�Z�pY�K/=�^��ڦ���h𪣠������CM��l�,�m���Oj�_�iZ�⦫��W9��?s\��SHZͣ�?LĖK�?*Y�os�St��{z{S�Q#Z�>�~j5���R��l�t�W�[z�<�Hé�A�H��q��^��)���u���X��My>���;�}����ƣ��H�jX*�A���(s�Ȩ˕��qk6��{U�uW���ҿ=��ڋR���7��]�� �6��ŋ����y�5-N�h�}̗�i>�63��#G��|�c���'<�kٴ]j�R��.|��2�c6
�5���n�=:K���EJ&�h�������1��M>G�۟7#��+.R��=۷�Q�����?8�y��چ�^������
�o9�v�E�z�SE�%�)<�ZB7�����ڄ(����jY���f�y���O^i�U�ҼR��Z�gvX���hA�-FE:c�6*�Q뱈���m��Z�F�|��W�A�mFn������H(��}h��E��N9���4l�-�3�^^5�On|� =�5^MwU�[�V,z��5=+ŞU֓"+n$`�k�����=�Wy�N�U[��G�����h>4��dV>Yn��(�#ڼ%ao=�yʍ�@�N:V����c�L}+#�WK���A���+NmV8���sZr�Ǆt�:ƹ�Ⲯ>�WRy�l�����@%�0wnEj[�*ۮ['�B]G}+�� g�kS���)\~��'�V�!l"�+�u>o#���Cy���{
�I����� ���)i�<?�1-�1��_&��឵�\I�I
�1�����k�� ����%c�ׁ�%��1Y#V$sZB��3�5#�FG��6�@C�8�E!��{��_F�^�.�%��]1��L�ץx����6��qc"ļ���^�9�#�J��d��@���s�|T;v�t;v�3��_8L� @#>���&m�{)��V�gu⋛����1h#��s������r20+�s���iٮ�67tqӊ�f̬�X*�  �*�_ �m�{�n�rI$S�c�I�s�_�2I�ʑ֨�͖������Ef��w�+|��@�Ŏy��l��42���Qґ�� ����K���}i���?��*5m�8���@�G���o�}4m\2޵�����^���ߗ;}�ҹ��waw6d� \N�z�Q�>� �^�����l�$u��wrT�=��1޸�H�h�1�99�re;֜q�c����Y��&�gץRԉ{��3� ��Tu�O��+!�Eܫ ��y��8�:ו��H�v��<t��F�y��k#�x�%؟֣E#C�v�����bkI)Y1�V��>ſ�q����	
�s�g�l��E<a���ú�]�Xq[SN�%i�+	�N;���'<u���� ��T�"�8a����n\�:Sp7g~*2�g��犇�ŉ�&:H�W�{R�͓���4�� d��o�=�Jz�?�1���=x�n
N?�0�)��֤eV!G#����2G�iv��(ʳ(� c?�J�d�Q�^�� ?
L���beU �=9�1����$~&�T�|ͻ�`���>g��րګ�G=>����N;�x���*`gҀ ����Xy��9�.c����x�	m�2�����'P�0���Q�6($�p;�Oo�H���h ���q�1�}=���ǒ3ɩ�(�Ԟ�� �1������8�Ul�q��� ^����{�K��I�v�ր$L��^�ߙr#�Ԍ������?�#�0�_qAC�j��H�5%Q�m��0�����U1�a��ӎ��"GG��u8�K�UH��4�ŗx��jX�� ��L�li�9��Ka�w�~�<�=�٨��U�?� ޼��֜͵���s����B�ۓ�P�S��
f�8���)у�8��#� �M�dhW!��Q�7��#4NÀ�3��5Pv�^x�(��\"Ɍ�
��*�_E��<����\����BpO���p�Qʮh�3�k��._����� Y-�z�}=��Y$�O�����3J�`��9��+ڳ�{�I�wZ��d�9��=~��H���ǌU��wW�U�4�OP*$�u4��u�����z��˸�s�e�?�z��>��_\���P��X�� �若/��s�՜d�ƏmNj�xx' �J��I%w���8�U먇��T�Np?�S�03���:q]H⒳)����NT�'9�;�p~���R��� �?�Q"���_�|�8��K`u��L�0z��H�M�{r� �Ui��a0�&�0�Ŕ��嵥��*� v�"�rc?1��H�31���c(f�*x�l���OZCVx�;�e�s]v��#b�dr�W 3�	Zj)g$}���:�G^�k��ڣ� �\Ґ$Ё׎Mi��mJt��e2�b҄�l�̳L�N��]��-	8�A��5�M�Aϰ���F�1��?�J ��^���k��a��]FD{�</j�g_6�9,q_i~��������hهs�q�?ڜo�"N�掛�?�c�	��m�!�P��,�")������ֳw��|3����[��h�,rz{�4�������цy5n�b(Ӝ��\��?��ZK��k柌?.|1rn"L�H� k�<��V�ҵW���U&��?�׿n���
(|�N�����Y�-Ơ�P��U}?�U匎O�,j0@����� :tJ��3Pnj��5b>b:V.�1[�1��[Q�*)�sڌ�k�z������*1<�s^���jo���>蔨T��������{�{z���#R�Ը���	�iMks~���
����_	`٧�����z$������W��L�K��i��l�H�b)�{7�K6 �Z����Πz��?�h���zW��0��YvaҖF��7�H����|D��B<��?�Z{��:g�+�-�����k���[�����< �Rw.(�I�]Y����Y�b�㸎�r�"�)���A�'�½���Y�T�9�%���͵�*U;��Y�>��n����֐��9�@��:S�)6�E '9ȥ��n�\���M�I�s~t|�8��y�'�9�l�`n�{�!y>Ƒ�^_Zg��RCs�)�$n�i�� 1�֞�hU
����Z�8��P2f��dU� -�¬�2H�i���I��4���Ѵ�@��t4Cm��N�]�����h��眊��k����q>�jk?AvF���a���94�})������b�\���|l�9��5۫u�o�:|����z�Gs�o�Wp �>^Y�����G�WV���?vn��,8���0x~�n>`�)l�ӌ����𱭄eT5���4�;ĩ-����C}��<�{B�D��*}5������L�<�jg���#w?�}�6�k�x��J�o���y��τ�U��$��շp@��B�c��F/B�Z���S�8�"�s�����4x�N�F{ud�Al�Q\� �M|�/����y
0;� W@�����Z�cwd\�o���V�q(�CS鏊Z>���K-�����
���^{��i�G:�������K�����om�A��M�dg�[�D�n���;*�����&*۟��ڥ����tehd�X�����s�m���`�H�T2�������~)G�&D�|���k�_ن�a�Y eY����%��՟������ɼe&y<�m�U�t����ה��+��bc�ק~ғ,�4WU�����ו�e��RN2?�gԸ���uh0N��Z��Z0�޺�;f��F+�(#�Yf�l~v0>�i�q3��#ƚ
���֮h�'`���ֳ�<�n�u�ѱ��zA$���"����"is\|Ѧ��!w�V���7�7J�XÃ�+�mA>eǂq^��A��� ���n������
�|>��V<�r����O��F�9�ҽb��펥��4,�� ؠzu暭�Z=�Y
܎��V2n����&��I2���_9xz��� �ۻ(?�k�� jkY#�����ū��'�6��Z�(�H��_��c�Y�U�>ڇ㖕a�����{�� �r76:t��I�> ����n�Xr�"��<p9��k���|��D\6	��ʳd��?�>���g ;�-��+&~�魶�q����[�Q$�w\qTl�1㌭\�`�ʑ�#��9��)-�1Fq�5v�܅��ܐ2h�����}�g�x����A
�c`g��^�x�����z���/1o�;61�=+hPѵ@ �61ϵz/��G���$�xq��yΟ1m�GN��?t	5�:AU8{��洝��4mfhY\s�ߖ}k�|?��H���A�8�t�8���ɘ[�"�<��i̪�{�;W���Ҥ��FM�@��3�Z��e��H����5���ۂ`ںKF<M�+�#�c�c}����u�r��^���KⴲmV���_ֹM��9T�F:��[z�֏s����W�� �Y�ܾf1�.�����C7��v�-����&��i+<k,�!}�|����m�	���ʊV-Y?*��F�dɕG��_�V���U��0Z�;y9� =���?���U�m+/��� �V��{[Y3%����������Gs�[_����$�n2+{M�ɧ\.f�p�?�|wk�I�}���?�kB�ė[6�n2r}� 
�����a��Ҷ�/�⧇↚˝�2>�5�L>$�܊c�9���mR$�C��j���Ū����4]N#�20pA�q��KR�4���,�]���+�#��H|�&�G�O2P�p���<��S;E{D{���R���4S�\� 	��5<?��U-!f���k���������Z��H۶mj�`���{���	{˵���� ��o�KJ#E��n<�z��+`�ǡ�_�ӧԮ6[��[��=h�"��і����{��'��i7�����G�b�V�-�N��ܫoS��Q���-�>�� *J��G����^1ԃ#
+��I��Z�/%�m�6F��5�m�N���ӭ5FHJ��k�~2��#b.uU��s��U���'�;�֩sa����19�q����_�o�������]���s�]w����S����VX����3~~�+ХOݻ9*�]��X�:�R1����Jd*y��kL��wexW��`g�'��Rĳ� s��Zס�-i/�Ka��x<��Z�w �qW��4`�W#�:� :�#+�0�g󤊱��8;�+{Kӣ��9Jd9�j�f��o�Z����kn�b�_�Q�RSG�ftn7(��U$��qV�Meo�ʏ� ��P��랴�~��t�W<}sI��y�4l< {��ԣ?t��w�TH�aU�2>���YZ�Qʲ�FQ��u��V��S�ߏ�HŔ�ۓ�5-hK��7Gn�l~�x%��˴�<����u�kϙJ�e�g�:�� ���*�l����aS�;0��)
>�EL�3�jI?�?1랝��H95�z��ne�<u�oe�ӳ�e��c���|� �����`/�̠�,��8���U~y�.㟛= c��vu9��b� t��Ē�J8l|ޙ�Fǈ1�m��x,8���;�������J d�� � {ոA��G�UU��Q���4j�h�5`}�	���8��/��6{���� �Sp�6��
b
�ds��s�֛�rH����}��N�cr�� d�O�|��e�?�h( ��� c�q��H~gs����.���9�֎x�4 3�s�tr37N3��g���J0 �4 nx�89�ݻ���Oc/cҞ��FO�����Y�:R��'$ds�^�cf�8�&H��N	n��Ҕ����'+��|��j���
` |���N3�s�)�ۛ���zUc�0<P���##����]�I9㨤���瀿ʕ~e ��uP�'?��\T���$�s�C���S֤����dw�� �m��9��,9U����Jr�H+��s�n�}ݧ^����0 n�� �� ק��:�����TxV�~W�� ���.� 8^�;sH�/#�֘�q��Jsey<�� 7^� ђ�}@�NўG>���X�����I�sL�!��i�9�a��/�� �SFr�)�Ԛr���6�;/���#�I#s����+'���ڧf��G�j5���@ n�O����\�'8���,m��������v�ڤ��hs��@=iG�����Ӗ]��t�Ԃdݝ�$��=>��x���]���0��?�&��]��q��sU��;a��
�c�Կx�����U�Yؑ�=�6���sHz�ݯ.b�?��m�/^�U�O¿������5�%�`<��~g8�'���_-iW���\ȹ��8����<e�i夑-�Qb�-�h��w<�ҹjA��$��~ ~ж��riz$1ƄV�����k���g�n�u��9#�Y�c8'����=*��|��rH{f��yN�.c
�2��$w��;���HBc���Y�E�ܷ��+l�H ���]q��Fdy�bz�)S�,����H�sc�Q��� m';j��[�\��?J$̨O�W��$���:��U�3��I�{K�$���Q�� �����t�)_�j5�:Ҝp�8��:�gw�1�|S䐳.�1�����~�ޅa��d���R[�A�=*kY����UL�GzO4��:�ʀ:�8o��]�3�ֹY��=��N6���]��o��=?���w�d/�<��`1�f����t�.���`J��⹏��3]7��m� J�<�mV-�wq���2� `A�˰��Ҿ#�]ڊ��N�s�_Y|�4;Y�S������g.���o�|`���<���]�s��־����mt]�A���W�>�..�%j�G&���r�?wq ���Z��w��s�����xu+��=�t9�y����{��6�Z:��FU}�Oҽc�%ǝ���I�yG98?�_4�5��N�� 3ɕF7~s_A|S����-���>S�� �W�K���\�G�q�UW>��'��4�bU��3뚎2[V��G�O��7oҐ=��	T��n1���#y�'>�5rU�9=�H�Y�> �t45�67\�������� k[(�Y����W��nbI��O<�?���������}+	ntS?F��� f�?&?Q]ԙ���\7�<6��F	�3v�����QWNG�\'�<T�M��>0���L!�vc�c9���*x��E�G�֩��è|Aֿ��yn�k�|2����)$Qq�Fy�|�o�@O�<y�z�u?�f��� �@�������e1H����s\'�+�i�x ��jw2k�H�1R�WО&�V�����vg��	|�V8O�z5��oo,(_��>�?�_����5ݠ>Y9�����:��u�+8��:��f�=cHp˿rJhN���s�&��[iI����T��Y��G�5�7�爷/ʻ� �{� ��A�h�9�Eַ7����(�R���i��!���B(�6�9�$��=9�{�#�I�ʊ�|̐�si��ȫ���@�0�<Q=��(h�z�P'�c�6�v�|ǚ�H�`�R�.7x�����cqc��+��q���(ٛ�]Ɩ���zb�?��Z۹D�M8]?���xu�n�
��5���ӡ ��'����,O^��\@�0 ���92}�M%��[E��1NfU]��ז�R��i6�>ހ��O���٤
W�k���������,"gL�6q�+(h��čx�x_��l`��L�W��'ផ���/���wT�6���mj@����~�/�}k����$�����,d�#eS��������z=����+|��Z�-�����WJ:�u;� ={�p��ֲ�]�I�p~;�ˁ���cSb��G�U��M�
-���_�oPm;�q�[`YO���~�|^��].�V �m�U� x��ϙ��\�s��j){�A��Ϯ�/�Ik�҉p�{F�\W	������$��\#1��<b�w��&E0���e�k28.كۣ��[ֵ�f
:X��㿏�<W���24�r����Oċ="cmtT|� ��ۋ�TF"����Tb���]��=���c����z���x�#�D����5��B��g��r��6[S_,��n�-�|��f�n���'�t���5Wd�X�[ԟXդ�nIc��{/����~����s��Mxxl6Э�|U���1�P}�o`�y���7��>&iW,���� ��63������&�V'ڵ-��ʧ=h�v��?��``V���mc����\*���!
����*��hU��4��徰�c�������Q&6��}ǚ�� ����Yz�#�;�|�����:{?�~^P�sֻO�d��do7Nz׏�?.�v�j[}]����t���g�� l�?K�%�� pwÊ�տj��_��8��#��ǃ�$�҆c�3S��Z��� ��YI����=;��ě/j
��	0z�N*���yg��R�a��v�׎���([�3�kCM�u��;�_1^?¡ۖɚ$��_�����;��&�rÑ��z
���Euo��2W-ߎH�W��"���-SK[	��`��a�}��Ξ"y.�q�MĎ+���ڜl���?洌z���u]�)#�Z�E�x°*�2E7V�d�;�k�&��'�Ky�E�zb�o"����\�q������L�w׏J�����ec�s���W����q�9�^!p�n%BK����oL�{�Cu����|[-�s²m��=�ȯ!X�\ϱkKզ�.C�$g���И�3ܵ��n%V�nr*�7"�N{
��"Eqn� ���H�V�񖞹Ċ�<��gB��k�����,X���l�mFw)#��;_��q"�9��]|P��d�~'���JH��ﯭs�85����/ n���L�9�����-�d��)��fU�e-ׯ&���p�����\�d;�^�}b�X�YV�#�q�d�~��;Z�ԾK����zdWo�]jWLcl��9�W51���=�O���q��� �U�� h��i�v9������d{�����-�3�'��������E�)`�?��SC�+@ݽ-�R:�ݚ���/pѰ>��Mm� ���Ge9'�qJ�,Ϡ�ŏ"�P7l?�'�F���ͤ�xϿC����$�����]�q���z�9�[w���^�s��Z��
$D��� \ҷ����������ϑm��� r99����Yrx�s��KM�}#g�o���(9�q����V����ŀ��Ռ�k�����Hs��q�j_0�����;4�-��ö�|�����f�����:�Y-_��݁��ɱ�nI�� ʥ�Cg,��K��m����7�O5�!���f�ߴG���n��R���k�Ʒ,ܗ=��R%��	l��������ϒ�~��0�ѺĤ��.3��k���U����j���^Y�G#'�֞��ƃ�Nxv����Xr[�W'�C���ִ�/G��i�c��H<���j��E��b:����1�0C6S����{Xe�8�o˕Uw�7j�2 ��	���D�.W UEw�ׯ'�{�`o�{$����d�F{����������.pv�s�v�� *��א̨~��Z��,f���``@4\����<�g��N�W� q�����,܆��#o9*����¬̓j�?/4�Jv��C�����Ə42��3�@w+��RZBd�@�< N9�W��e��R��5�.�.Fh��+�\4R.�ۥ!;�6N*6�n�n?*�Y�0�OL��Er��<�-2�����&A��n��z/ʸ��?sp
F::�<e-�.��s�i��x�����{)��=���⥃�>�ۓ 3��>��zD�۳���5��`K��r�H�G���ʽ=9�z�����Р���n����U5�G��f6���?��3�;�8��������ڢ��7-ic� �z��G���cn��B4����Z�_O����3����*��S�A��d0
�@=�֭� �J����j� �"�y}q�=zv����{[(�=H���E�S�X�>��3�[��ZKᛘ���q��K��p��+�9�c�4���َ�\g� �J��8�L�� �]=��~���zc���Vl�!�pw(<�8�3G8��3Y�W׭2C܎:���K3csm�w�M���`Y�E_2#��7����P�d��)|�\�]����q�S�
�0=zc�QF2rG�H�ۈ'����IN�� 9v韥6O��S��g��I����3�Ӹ��ɠr{��� ����y4�P nݾ��N�ހq�WsޥYS��7r�Am�M9��$����Ҁ���օPT�
�c(!�O��B��{PdP�/_cȧI0*�W4�b�	�N;T�jT_�(A�G9���!��>��N����0M'�v�z/AӨ��a�B����,��Dś��)�z���S��*Ó�a�ֺu=@d2n�����l��s���y��3����5���Z�:!�o(�����N��S��
?E��0�]�2w>2H�S�|ʤu�[P�p��s��ڬ�h�M�![�K�~���3�`2� Z�4w�&�I�?m���Iϗ�y�SG��2�(����O�ٜ��� d�d��J��%s�(?�vv��V$�P#���j��=�B�(�3Ȩu�h�8E�0�i�)��d�Skdt���K�R*c�횙��5�l8���}�s����y�Z�#/��'U�>�i�nŀ
�s��zLpY#��y���@��L�B���v�=�>��}���Nz������F�T�`c�����i$���3*��Gz\���s��le�RT���Qgܞ����)^�8̊s��n��>]�c#'��sH^�=�<:M� ؒ2s�aҮw ����{��{;R����+�;�1�~5����;Q�!\`��=�O�ú��to�֮��y#�I$R n�� ��n������N�҃�M�pw~)�6
#�X��
[���Q��>����o�H5(��Xg��W�#&7
1�J�Vktb�X�@��B�\g#8$������q�I#�k>ku`H`>��5�|�)�a\����՗�'ִ��[*Oɧ��6�����12g�n��髀�FI��������b
�Q`1��� �>f�G��V��M�ۆ��n-�_�nX�o� �r U�#�c���>���C[�.Kw�5E�+�y����7#&�X�#8�9�#n7�jз�&L����
��i#|����L�6c����M%�[g88�z�fR����� �7� 5�hr�
�dW;�b1Һ|��Nx�c.�n���v2;s_Q| �G�US��.��o־Z�SowܒS_V|G��-U7T �rW��[��-'k3�ޙ�|D����oC�������R�Kf
��_0�\]x�eԒ����*rr1���5���$�]a0w}>��K��w,G,O�|Q����_y�
HNs�{����9X�c���/ּ3�W�-��������\q�� ��*�_�P���MA�$g<��+ЧXX��4χm�,l��)[�pA�I�Eb�f�iv�=;�Ԋ�VU�+:Eq��ѻ�A���s`���jA^�^.y������ ��ł|���I8a�x⾎�/����y�>�V/s���;�I�yX�=�����?�p� 	�y�����w2(V��ҷ[�,c�)S�<}+��j|i7�g��Wؾ(���&Noj�']�E׌ �N���w'���|΃Ɵ��44�M�|�6׉i>'��:��M��pZ��s����.�l��^!q���5�Io��Ƞ.�dl��GI�,�'�	?�{&��r�/G�K2��zW��Z.�$C�;}jY�.G��ġ8�	���Z]Sč2gf�+�=V�J]�v�5�_>�æ���?�l�״G
Y��b�X�K���������\�⻯�3��v�q.�M@l!��k��Cba�՘,*li+r���V=��e���8c��Iǩ�@�y��)���R�Z�לR){��s� 
���5��o���ұ<M��9Hmn����
3��6���ܕ��89�='P[laj/0]�e{� ������W���i.wı�=�ҽbht�/\s^i�F��V�6���4ķ9-×�nY#Ry�h�,%��B�ɮ@��Ͷ�&��m5���<

cu��&���k�/�M�j�$o�_G�ډ���\uǄ��S\4a�}�(l����6����g�2��n��k���mgR��ӡuL�x�^�}����w���^1���>izj�aRG|PR���f���d�np)��ߋ��"�1�3_gG�=.��?*�o��U�ނ2;|��W?�����+�0ȱ^+�W��_ŋ�[���+'T�7�N���R^�
<?��������b��F��+���� s����6�ן|S�ɱ���aSb���g��M����x=��;�Lw3�~b�����Gt� �E|�y�H��95��.�^�}ϊ� J�L�ǽ}G�o�v�ج�[�ORk�k�Տ�pL�k����V_�Z[/��|��G���wB�.��|U��n���u�U�g[K�C��z�ß/5���,N����o�4�k$F�s�y�XNrZ���-oٺԞ�>���~�0G	XT�w�l_�cq�.W�x�� ���
�Ҡ�������|�߳�������oi� wG�D��\u�phq/�B{z�o�EI��O��\�����L1�>OS�K/��m�O?���o�z9���4�����@ލ�CS�%ܮ_#�b��Z+��C�;Wq�| �Kh�h~U���v�|[�#�=2{SW������(u'�9Y�\��Y2x��G�J�c
c�Z�$�ǧ����Q� ��Ӄm���=����m�|�~Q�ҡ��9s�_�95�7,Y���O5Vo��r�(R;����S� �d��c�C4mq'���k���r�Z����|^��l� ����-?��?�s7�����/Cy��a�eET����������f����rܱ=�S�>.Z���
�� J\�B�f����?PQ�%���)�xR*��n�zW���~8��b����a7p8��J��}ϰ������r�)� ��CĜ�@������g�oʠo�N��s0�Gٷ_ nL��Ro�E��q_/ũ$��M��d��bO֗4����R� V�Z�%x�ӽx���u(�De�	��^�v��q������׊]e��Ld�|�������n�������aU1���d�W<�<�R[�<�����м:����C��<j���&����vF�	�u�X.�upz|�z�*����bc�=���ⶍ�OJ_/��M5I~p8��y�x#�\R���n�� :n>\���O0�>h8�z�������[<^����9�pTd��?��W���.�8�]� Û�]���7j�{@��\�Cl�G�G��dF��T�x��-�0$�q�z�͎�pV�};V�C�E�c�G�]W��K�W�`8�sڼ�;��� �+��V��hX+�z�S�� :�5f?ⶇgo��YDJ7ɴ<�	��?�x��Ķn�~`�r0E{ĭU$�l�!H�R����^-vVi_x�:��uR��d��J8x�r>e�:zפx�ͯ�!w�wl3d��㯵y�w&9�<�zf��᧋�lt� �Q;3���rzh(�ަ���;-b[]ϵFW'r>�wO�1.�x��ّ� �>�z� Ķ�x��d�e���6FrO��V�7���$�2�ޥ�蠏ι�v7I�+�]�ýR���,��wU����qSB�$���W��ƃ>���,B�6�RM.��,	��~u�Mۻ��(Pzr=MmK�1����:�L_1d!���V�}Yt摤F���
��}�ڪ,�fgfR��h�5���!R?��Jz��@�*e$簦��F �p=1@iX,Ge9 R3�d�x�ߴ�#��=0F>��i��N�3t'���f8l��/�����t^I��8�jl��42H�#!���ƣ�M�]�UF�`@���fx�$�~��u W��;����A�k>��c�L�vW�^�P���rZ�2��
�ҭ�R$��gkd��Bj�'��v�Q�1V��#Y�>���)~��H����1��A�'�x����~��&����*���Wd�lԍǕ��0z���Z�V�r2$P}�1B�\r��8�\��VZ���Eic����z񚴗Vq�O-\�G�ӧ����ہ9I��Lα���ך�CH�=R�5UPc�E9�ȃ��9�לy�/��9�,��2u
�f_�g�6�nI��R[붲�$q�Ny�6G�I;�?�]J��Əf?n�J�Y�����@,?�/�!UQ�s�y�rHc#q�|Ő�_cu�<� J�f/o#�c�]��gc���Ն�%���3/�0�~n���^o� ��1��R:��՘7}�
~�=�=�^XLr�3|���ҷ���p��sXr};q\3I#C��j����`��ϵ?f/l��?Z�9��n�=>���ĩ"�Wۓ��p��/�X�\�@;9�}3G��gt�!X���z����*���e��ٚB~n1ǵ,{��l�`y��Y�Z�vK���?�X08�5�Hdc�;��?�(8��ߎW*#�]��o������ҳn5&�b	�8���o4�뒿ҝ���rx��C�f�_�]��q���>��7�U��� xb�$ʮA��Dd�!x�U
��`s���T�d}��O�e-�
kq�����c�C

��Oj<�U;X�H�9�ҝ�?)�r.y���\R�Ly�9<�I��3��ą����4}&�7�y�*�j
U���b�Y����w|��Ґ^�dl�Ü�ґ���?TZN��Tq���Ldۈ��J�#kyFl{��p�ri[�|�Zr�7�Uwʽ[�'�}����i-������iW+��z�,���@������'�`a����x��I������\ӓ�Wa��8�6�4������Ƅ�=G^)�X���+�m��i*U�jO�W>[��r9�Y����ۑ۶z�d>f^�ظV'�h�?�9� �Sd�'��b?(�?^�j��~���n��ڝ���{�r����͹�oӽDu��d|�����sޠ��8�~�Z6�́�����A�"�k�;~���z�m��.p�rz��1	ܤ���9z�z�zqK���%}j�~2�(�Z�U*f�:94У��G�C��qߎ�X�g�r��-� -��$��̜3�})� ��#E��9��|ϸ�\�����Cmf�j_![#�֙����E�6b��D�=:g�=)[S��M�3;���< E?�i~\�G8�ދ�G��|��G�2��� a620<R;���Q`!i�ݻ�����ҕ.'\�o3=wg���4�ʹ�t�D.�2�7����MV�?���jv�A?��ن��H�6Yc��O͕�
�N���<������� ֪��2�j��J�N8�V^Oܐ 
ERo�q^,\H�!�親���$���֝���=Oz���8���ZWZW��Jq�:��F޸�H�Jj�T�=�i(c��j�x���^zU�^�I
�M���{`n4ؔ�\� �Xw�	nLm��+B7����d���U'+�sC pW �GQ�t^�l|`Ls\�*��Z���(���z � {�bp��ھ����]g�;��3��rNGO�5��n�����z���,�	R�Z�˕⥡�o��X��o�[�k#�~&�-�L��d;@��zׇh���,�;c��g��n��}zќ�#� =kU$g��G��G�L~���U�/?6=~��~�_,t��ټRO0�Udh#⼇ğ�&��ۘ�?r��ʣ?�+ȵ-J�_��]��+;|�߭K���#M��r%_*�I����L��� =�i�igj�s��&���P6T���I���S�A��֯�FUI`�O�y��^FI��KgØi;dw�}�Q��Ű�h#>���^�y�.I��7��j;�����&�{�T�?H���@q�q�z� �k��s5p�	e?� 7���Z�xf��1#�E��Ќ���~ h�Hמ��}+����_��Mv�Y�O�d�1L�����uO�;�qw�3����5�%����t���÷���o�c��4��@[�c��\-�D#w���~�ǳ��/�_Ӷ+�h�h&ID`�ӊ�0������:U!-ecK��&��0�1��|Q���c/�5�?�y�q$v��񗍟Z���św -2y}�LmB�Ox�b��O�_Bx_K]+H�q��+�~���K���'#p�W�� (���T���i(��hrǩ�)qג~���z^( �p:]�S��q�kc�4 ����W;p�Ҷ�����3rAh����u���p��RH�[�-�O���q].�n�pȤ�wZ�-��r�К.՜�e����7�|%&y�9�z+��{�����-���pRV�Б/�����L���z�h�ڠ^��+����t��+Ҵ� :�3ގ�f�҈S'�e^j�D�3R���z{<y��{U�;�}�;�9���*7��x<Wo������\���Ϻ�_��Ͷfc���q�|L��YK���KP�����E����� �d������@x�=:S?�z��6�G9��^͟V��k[qî�SOG{'
�W�W���~m��wt潃���;f�%G\z��c�-\H3�+˾2\t��pq^�
��Q�y?ƥI���ұ��T�$~w|Z��mB�1���^s!�W�*2zW��O]ڕ�|f�J�έ�	����g���"�t���.�Mf�d�z�m(l�@��	� �W�iZ��,��B�9#=kZ�ō�Fع��g������O	��C�x#���=������o�~ x��p�p7}k�� ����1�)]��Q>c����0xf� �b��T�7x������&�]�ً�j�j^�;�2���m�|��[�P�~�njp���k�V��ݕZ5ʏJ�ɳ�;���|�/���%��M7�z��0����춒FF���њ��k{
�q�N��g�M������e���9<{�aݻ�5�T��W6�0 {���!�V,����<?]�	 8=����K�?:7���{ǙkU}z*9$�T�q�=��>��E�x��YK0'��r|9�����kۭ�m��ð� Z�mJ�$	� O�}�E�����|>�T�cm޴�|7�hK`��5�q�8� �s�4��-ռ��?x�􃝞�n#�v�os����{�Ie��@�Re�x򈣱��2C�#��� 9�y�3<9~N��O5o��ȅ���+����i�v=)��Dc#
W�j�	�<E~͹�����|:�TiQ�ׯ�*��MjX�iuj��㡥��x����Fu-�V����
<�9�<W��<*8=���l2.�v|s�&s� ��n��^5 V�V/�'��9� �W���� |���&�Z��s�z�ֽ�2�@g��קЌR���*l_}������L��R �{����� ��g���m�*{��T~..|X~a��q�l���?
�r���M�?*�s�q��Ǎ��u�g}�����C��\���q��F���5n��H�©+�4�����N�;b����cO�4�a�O��n��6��94}�7^v���֠~7w9=�SK���0V��g>޿��t�x����j�� ��ۛA�y�K��ݶ�� Ҙ�"��A �y��K�s��&Q��@]����xf�\1����D����8_|d��8��Z�����S �5O�ݖv�(�c�Sn48��x��q�d~4ְ�3���<�YH�Q&��K�iQfB�15��h]���1Z�R���z��-<���<�j�˰6s�����u�V#k��ʍ��'z��4v��O֮Z�ok'��}q֋��_¬�dE<��V�_j��[�I�%S�O5����E�q�pj��3 ˻pɣ�4./�-[\��:������.�p����\f��%���\$aGlgҴ|E���£|�x�ޱ$V�L7O��G-�AqTT��,e$d�s���iW*�A�y9����B���1�9�)��oR\"�H�C�V��<9g�xH�IQ��7��mL�\ջn�F� H�F��5�I���H��P0 � C5t	��P���BC� �׿#���*�T��A�;�[z/�.t=6�+s����Xv�J�*�Kv�'�N�J�#��ν}{Ug#��$g=x�R0S�w�⩲����#�~Y�����<���~u.���>W �S�Y�ut�� ���)��@�K�k�[P�^L�I8�x�������&W�$?t��<d�U��x�{V��+m�0܏Zə�s|���������B{�`pH�}qI���>�GZ`�ʹ8?B8���C��Ҩ�ʸ�g4��	��'��M�rrG|f��=;��0���=qG��z(�6�(�8�Aʓ���)I�
��)9�8��C2��A�zI2ˁ׽��$dP �V�oniN1�9��ʐ7Ĝ�T��p� t�onhR�q���N���)���(H،��� ���JX��)$S��h e��ygw#���n�ޣ۽ /����R~��ߚVP[ �;�SX��M��5�nr{�C(^wå1HU��h$s0f㯽.�)�n#���,j�0
�����Cn^3�<Pr��dc�ZƎ�L����Ϧ?Ƴ���p9��H��by�z~�2�^��A�TA������'�R���h�>^X.��B��s���wˁ�(�Tm?)�� ��A����1�N2q�ME b��v����w�*OjsmF 1�V%�������:����5�S�ҙV$6ё��/����2h� �_=)2����҆��	)����?Ŏ��21?)�=8��#����8���j�)�&���@c�����X���s ���@��N2 �&��o z�|z��
�7��	�eS�>�q�>R}jnp0=��f���Hd���i�B���ӥ7w~���-�W�t���0T1Ӛ�w\����S�9���A�{��]�>�S�#7˜��� �L���j9*;���ջ����Y�¹�j5Q�c��Ҝ�۞�r�n�Z7��zf��7�=�\�Gӡ�!w���7qP���Azz���.� *�e=�\�ךQ'Q�tɤ� |�sC|�B�����*�ۇ��H�-��֚�{ߊS�Zc��Mߵz~m<u��t��U���sC1�e��vW����|��J�f�x��N-����"�~�Ъޣ�����^NlR. ���T�s�N٤�['�z c��=y��1&� 9"���������!m��I� �0�g���Z�EW��L���H��:�*JU��~���*��N
9�Q���Ѝ�j�Fx�*��#�y|���jhذ��q�T#� ~���v������a.���C��OSں�V�x�Jb/i�X��"�'n��u��<�cK��"�csw8?:�	��u���I�Ҿ�����b��=�玿�5����<�o��	�D�{�TV���LJ��(��+�mẐ�
ݱ�%�=�@'�����V�O�W�y�J����8���Y��i�i�Y-�.;�vrY�w��rk��x�A�҄Z���ǒ�+��;�_̦�Z�?������ ���`������"ƻ��rp+��(G����6�l�d�zs|�~󜑑ߠ}k���du<WD/k�*�v+\H&�@;Jᇭd󴃐ݛ<֥҅��&��R�J�q�֌���2� �>�9��3����}�+�O��h�ݹ]ų���}�\� ��������꧱�A��S����»����~��bw�J��N�;V�c�x��8�����iU�PqH����7:�ꢹ}�7�=�Q�nk�o���� B@���Z��OZX�#(f��A�;}3tv�������5}5� �+�� ��n�(�2[4-��T
��H���L
yn½_���ţ�����SZ�������[����Xt"�NNZ������Q�Qm�sN�/�zqH&�d���H��h�<+�|蕾�@�M���7P�p3��F�h�x�U�x��#eXS�|����U/$�IǽN����R�]����˯G�<ʷ��Hܶ�k��=��Ï�M�H��]Ž�ǖ��9杀�I~�I�+�<q��&��<v�R�O�ie��y/�-mIUwa7��Q����R�F
zu�d����)�1^K��.-UO��9럭{%������ݯ��4�,�8ʰ�J����n�����d�ȯ�׷5��h0k���f�EM������6�K����Pp����C�'���cmõyo�σ��u%ͤ{t�+��� ��� �!�\��sO�ѫ�j��ar�HW��Ѿ�Y���Ms�����)��9�L��x��Ю9��C;˫/h��tL2ġ�m��S Ux�>��Y�m�4$r�ּ��S�{�=�V��t�+����"����V5
��~t�H�Yo.�)�$g��n5ˢ��;3m�f��E�-�����&�ͼF�ʪIb�a׎?Z�;�&�x� ������t`��J����C	>���>,ɦţ��P0C�W��W�)\�����KH�У�Ke�<�^E}���g�������bI3��N*E��BG=3NQS�qn:kY|x�����wzY��<�Ԯ3o e#����o���SȠu��~!�@I	a��\ӧmM�;��q�4�3�j#��E+� z�V~�2�Z�a����M�_��ڰ6Ca��c��Nj5�ES�s�59Q���:��LV�ub�����G���eìy=�Y�m#�=@��k���5/����n?���
��O�5eg�В9$�𧰬oG���q�x�j	�$����0j�H1�9=�5f^A�}qJ�-Z�*�-�s��ԭ!�s�n*�U'9��I�EX��������DpqT���5!r�����_��
��&���@�S>A'���Y.�,��(��KRv1���F�63K��9�Q`7m������@�e�b�O��h�03�>f�r�3�h��h�&P�gR�A��8��{�j�<�)e$׬Gh.�T$'�׊����>���i��7/�ҽŜ.�<O�N���7��M^���&�%�E�ŵU��� ^��9��WKmB�4��x��?Z��v�ao�_I�����w��iK�㾧�hk?���4d6q������I^p��mR\)�3����@�G𽘸�Ѥ�6����5E�[ȳ.���8��}�[��I3�[XհG׭2�K��2	�����`6G'��jxTɷ
Gc��ns���S���@�ۭVVx�3Q��9�H��*$'���p]E�o�ӑM�M˒TN�f���$18$t� �U��Oo7ӊϴ�xoc��F��B=��w�ii��N��>�'����?�����0�j:�Xm�
xc!�}N1�ߏ����t�>�LIIհ}0�?�z_���^=��H�.ȭ���7#wN÷J�n��e�|٪^}�HX �q�>O�G#�E��);�SҺ�k��\l�s�We���Q���%�FC�����\��I�x�!~�#�=�*�XdP~E ��־��� d�BM-�+���(ղ�����U��w[�:��8�|q�Ͱ��s��pH.��p����I"�v���'��_��@������ɥ�5�J~bF3�Gֵ$M�x鞕r����Vf a�=�c�6;x��z��8�*vX�Bv�(�ˉ����'����[RR��,�e��{{WW�*�� N9�n��1� hpwnʩ��SSp88~{b��r3�99�����)*�7 ���~_�[&� p�� JnI&�I�e$g���j�s�� �^�߳��l�#<x^�#�Rz~j��栤����1�����+��D�!�����,�*���{�����2����2?�Z��?f�iL�7�����Q�pQ<�c�����V,t+�JwXԻ�jZmևv`�F�ձ�~����A���J�d�H'�wG!��vm5L�G�\���$c�z݆ݡ���m���S�k�^ �^qTV+����q<�f�q 9�򾇟ʢ�C��T|͞NMc����}�_µ�,��p7qYN��U�zV�ؙn;��(��7����sI���֨����B����4�N��'O�ހ�7d�C61����P}M08<s��>�v��pOb:��6���w�ʃ���<����#&[����$m>�����w~E!���9�� �ߝ G���8��[s`����N�����ր.��g��<�N>��[;�4��Q�u�p���S�n#�(#�׵7w���۞�>ƚ9n�w�Ґm����޴ �y�Fy
phۜw�;l'<P������H7��#�� �h�WVۃ�Lb����sɤnX`��P�SW�R�(�a'���}��������=�w�N�?�ލ@06��z��B�ی�)NUN@�P�u�:t��ccړ~#9��r1�zv�L`T��u�, 3c9�7%�P�=��Ln��� h��8�j���rq�ɦ4�*�N��(j�Dј�`r1�G^�
�r��+�GQWU��CUf��G�p)UY���OJH��J���7�{�~(O����
���y� <R������)���H94tj�9�ɡ�ς���M�@��8�GN=�*����:�R�0 A�(i^��J1�c�4�nѴ
��#%H�ޙ�����*Aɩ2�]��P�̓�6z��>cC}���րhU�G��^x杜�E#7S��ژ	ϥۓ�)7u�v��@r�`㷽)��ҍ�1��g�Mr�8�v�uS��9�f��ӭ9_����۹�h�s��^ǌQLB�@'�ӾU�>������XB��#<���ʹ�J��֌S����Ҝ�8��F0��0�i ��i�s�,������n �+n� i�Y��#�ޜɎ�;
z6޼�`F�FKw�p�������������8�M�E��>���g�O�������O����4��k7����ҝ§\�b���q��H��Hw��֓i s�U_�>���l�}�P�6�w q�R�)	�<��/$����ր!e
�T���h��>r9'�s��P��ê���@��f�+�r1?*~���u��>�i^4��ɯ�~��۫�p�{��`��}}i�[Ya�x� m^��W���}g�ˈ�{+G����?h��W���+��Ǐc_� �A�L����4njEv�Ñ����s��J=��$���ǔ�����V'�ǥ>�ĚU��+Ct���2?Nk�4ԯ��}�Do����׼�ݿ�8q�z����Ƴm�����T��?����Ey��L�����.|��M����Y&����\�/��׋*j��OJ5=�y��Ȅ�ǽfɆv��Z�/� ��Y-�1��Ȩ4GA�4� �?�+菃;?�����5��� Jެ3�#�+迂�ͭېpb���M3�����8©�6w:�o�jWGS�x �U��[�oJ�ld*�^��3z(Q�=iz‱��L� d���GҼV�N���dv����z�!�n�c�W�-�Q��#���ۿV(x�O����Q2w�k6ŭo�Dy���G���G5�pF<�e��Z�J].�i3�"���U_Р'�)�z�4�Bq�q�W�x6����[4���k��m��q��*���^�6V�NFG�/Լ{5��F��J��:-N�:W8� tۙ7��ϾEV���c7��a�-��H��X�#y'ܚ�S�v���bEl�s⇅��i"�(�&��� �NÍ�k�e��� L��|Z��;�c��߄_t��*7��\�k���])��|��;z����iuK��߽{n�w���Z�7N��ѼR�"��`6zw���0?�OGh%�^��z��$!�-������U5+u��a84!���mt��*���U�8���}�*��fb��W�?�$3n9��.��0a��8�O\�9U�.I��eY v����q!VQ�"Q�i���s R
�4��>5�K�����W��㷏
�4u�M�db��o�s�o4�ܱ�|Հ��.�P��������τ:v�K��ނ���2��֬n<�԰<R��,Q8hHS�[Z�Y��2?ϭz\�j��b��	9V���ejmcÞENO�N�ߍ77J>����7����� *��~�y/�� �-�8Ⱘ\w?=�!�4WW@75��/�Tzf�č�D�������>����k���n�W��$�F>���-˶���M�u�����q��}E|�5�k;`���׻x���c�:��!�2YG�|� q���ߕ�fA�(�1K�贛�&t��t��S\Γo��V�������m����?�f��ŮO@:�oY�����2J��+*��Hn{^���U8�<�r�@S��Yv+�۠��t��Ň���R.��#��ؽ��E�I[O�q���+�g_���.:��!��8'�Qb��~"������q"l� �{Z��~K{�"���ORj�A�W�+m_��5���jKp t��ϋV+���X�'�c�G$ª
�|����-�x�s[�nYp95�~���ϭz-�e@�橮P4mC,���۾ka�VP3��Y�9nI�⯆;���@CMc��Z��sAn��q���=)VC�~T��
L�n�ңn��^6��8��
 :�Үm�	��ym�Z`=d#���0�; �j�9�Z8��M䖪dB~Nx���O�-���������v����}�r�M�@�\�s��%��m2�	���QY�r[>�ֽTqIY���]g�����{kC�"�F ��+����>]wZ�Ke�;K#�W��烞�_F�hZ�`o�X�J��:�G�^�e���Sd���#����S(�\H��c��~��%g�5�����>�[�+�e8�L�Z����ش��w#񩵍P*�����o�e��gr�X����rk^�W*�I`����I���a�6���}k	�%� �ӥn��:鯢���q��}\�B�'�
8����I�")���V�uYb`Kd��>��#�_-���u�ֲ.�\�3���k�p�q�����A�F߆A�2�������ҳ>�V�p� >��n,�F����5���c;��j����5�Ž����1�W����:����63IGҼ>9I��ӯJ��$d�eYJm�)��%5cH˔���_n<U�ٴ��[{ia���rk�9-㵹��m�-�S��V\z��Q������r�FN�U��TB� ��k�FY_�'$V�����+��� Z̶�D����_��^m������H3<Af,�Ȼ��qX����)�"��M|.��;�Z�bl�v�=���������� <��t�^4���c�\s��o�7io���9�I�)��Y7D�W�sJCF���ފ�J�
9>���I���4K]�2y�����@�C~U�KL�|э���rs�5�}��)o%Ď+�:t Z�y�#&{���f�x�E_n*���K}���h����M�eb{�]G�m�n�>ZI!^XGֲi#x��z�~-<O��������M�5��c�IP��dd��\��t�}^[#m�j3!U|����X5���r�yfC��*�S� �֢���4�Rՙ����X��)�� $�@��!���H5�>�D�e��f�� wd���}��NB��uf��+}��$}8�7�u�:��e�X�n�����ֺav��G�;=b��=�1��/�O_�+=w��7��H� s�sW5��͡�e�����c{���_���2�,O�ߍ���@�/QeR�#$��[�N9���D�qӞ���Ўs[Gbe���=�V��f�[�F>��Ê�E_�#�zQ�'4��u�9�(�4 ���� d�A��� ��y����)v�-0�h�s� =h�c?� ��-�I���~4�ғ$}�?�V�ӳ�8��L(�Dm���3�'�$R�p0y�b���2iP�|� �u%��i1�<��R7瞔���^�v�0)���;p-�����wA�j A�w�w�-���(�8�2��~n� Jd�ʹ��JF���9�g��S�� �����F�!���"�=OS�b�X���s��'�M�7v�`.q�0�қ��I�֜\�����&<q���i ��)�p��������
x� �>��z��s���;��;O5*N�����a���(`͎�1����p2��L�pî1ӭ"�X�c� {Hw�q���S���9�c��-�41�s�:���R.ܟJ3��z�F_��p=:��,rO�>���
w>���vp2}��ey�;��J[���⌖\}q�Sy<w� �O�_��!pkGL���9F��-�Vxo�6>�l��b���}{�5#�Pv��}O>�f��1?�^*@E`�iʣ�r~�m��)�������c'��0,��OlҴgp9�pi
��v�@[!:�=sҐ��2[#�?J9�������H۸>��I�)O� s�9���3zu�����I��3�}~� �^F��1Nf�?�5���4jH�_LR7ʹ�&��I��s�� ��I�v4�B�O4��n;})�F]�ԛ6�Fq�M.�pOZ M�F3M�^���7a�Ҁ�n�I<����pM/���q@�Ux��~����4��|gݤ�+>3��G�p'�p*ù4�o'$���]�4��F1����3��)��� #�Y�qJ�3 N>�69�R2�;q�LV�R>��n��z�S�;��r6ȽҐ�.��kwE��S�0:�ְ�Gc��4e2�1��#� z����/�T��pH�3ֽ��\~g�#|�=�x���!j�㎸?�5��W�1�ۛ�OҾ�+�����`qR�Aj+u��ҧ�2z���9Ԯ빔־���e�=q��ξ|���`ds�
�π�l�� ����[��TV��|f�C�=D���9� ����x��̠�L���xS��
���q�������Xg���_�2K�\ʹ�Y����|��UC�c�*Sp#n+E��t}:V���Ȼ�{VT��%H�s3�_���8�����W�?�=h�=;���Ze<�#�k��x]j�!��}{�R��~�|'��~��GO�滖�b;��m�����»v��ۡ�m�z�ʓwZ]�����Fw�a3iο�^��7kH�v�ßLWВƳ)V�ߵq��i�wɪL�r�6v���|I1��n-⑉f�{���t��@���$��gp9�L404�f�d�>[#��z�Ǻ/����vv��#�gֵ�㧽0�fx�5�æDN�Z�^՗M�|��v�ǌ.u;綵%��>ZBZ���?ŀ<ȑ�����#ԼM�,���7�� �/�I�_>KrwV�͠������4�>W���Ɨ>��)K�5�wĈu�5�2��c�p�:V����w¹{�.���^dL�(C�6��`������� ��?:���`�cG�^E��V��ȣ��kڡ�%���c�"DP�~�u� �kEW���Z�$�FNH� h�j����[���?:�3�o)��3L�R��v�Ƞ,z�s��;z�1�kk�H��z��s���9�7ō�s̞�I!��Y���h���*ּۗ��A����32E�νG«���1�4!��sc5��qt{&ϥm*��y��߮Kc��mm�RJw'wbƃ�:�R՚�e]��#9�H����D��|��|��L�\�翕�-) zq�kپ,khZ��T�J��Ġ���v��;��K�� ���6:��!(�Os_/�C��_5��˒ҫ��P= �J��|�|;� ��v=�ue���>���R��#֞��מ��� �t�N���
�YW{�3��5�� ��û�i�W�v�k��6�4k�yZ���Q�����ؿ�<��[��l��Q����+����u+�O�?1\�ß��|A����׭e�.��O��6x���·������h�����?�$l�y��X���J�TҦ
���6�&�MI��%��MgN<��H�m�J����zG��#6��w�y�����>:�S�Al�!A8��i3��k���Ƿ�v��Ɣ��ץxI�衑Tw�{?�~��ż��j��.{c�r7#ud���#�3n|����o��zk�|����ZE���������9�p�X�i$TW6�q��\3�s��K�s�i��V%��������W�8Ձg z�����-�e.��Ա����j(.<9s�+q"�qץ~v�V���\���B����¾��6��N��q_2|V�c�VRw)�?�\�<����\� �j������nd�v���5��0���{>��ïN�u	Fլ{T���[�x>�Jͺ������Ed2W�Tv �7)\
$mߑ8���X�9����1��X���=i���� K��Tr0��B���P��#Iz��厔�Gz �[�J�N��B���9�b��t�����6P�'�Z�� ��5��I�\ȓ�>YN6s���(KT���>�f�O�𾛢�v�mKPkX��`�GNk֊�<�K[#�7�W�waQ�F)�����_9���v�������8�������AЯ�Ge���� 7-� ����Q�]BB=Ҵ�T3��qק>�2]�#��-q��ǀ��\z��;�V�@?��5��1�\��=_O�Z:��lθ9����Ɗ:\�?,����*�Фd���sѱ�.��ڶ��Q��+�I�ҸK�	l.~e+�ڮ&l�I�=}*F�ܨ$�)�S����ӌaz/U���E'.���ZVW�o�?3r�O�T��'���=E$�U�p~b���m�h�Ñ�'��[�~-ۭbC2���0��x���占�c�����e�Q��8���_�	��#1���oL���b��U[���P0Ye�!A OqR۶�Ď���Vݽ�An�0ĂO�a���T��������"}��|}h����(�|ǏƳ|rzg���bܰ#=(^�O�H�r��z{UIp�yd 1�� ]T��-��=;՘Q�`T��g<�=(�����׀���*��=PJ����%��I�4�ޓ�� z�z�<3�[5h�_�V����Ҳ�*;�揤���<�8b �s�oj�U��V�������q�[9�y���c��V"�AX�}
��4��ˉ�ȍ�Dge��_9�~U��6ga�ˏҽ3�Λ'��YmIV���^���mx����ݻW�Z�&��`�ѱS�3D��n\jX�2��D�����~���]ZK��ۗ������O<��ǽC��g�5�Uu��&#j9��ڽ'�����(�m�v���z�J��煼	࿳8�\�m�����Xƚ��כ�����ѡ����v�F���J�q���?�]O��+��#2;C��8?���?jωx�D�7Cl������+�>�?
��f��;eq���_��kzi��V�:O]ٶ���Ш]�s�ֹ}R=��?(��jqt�g2�*5�\�Fy�R��Һ���!��T�fM�]Q��!��=q�Ù�H6�m�Emkcf`N�����w�5�v����*za;x'�8�F����Hg���8�?�>ԣ�z�n3�8��@U��z���x�R���@V�x��}E4���S�� '%OR��z�J�S��Θ
s�=iC������6��X���jF_��wm$rzR�70=h��ߥ(�wl��7P;v� �OZ.�2=��Fߕ��i��}i����9���bqNU�C�SY�i �:��P�+cׯ���, ʔ��րϦE7%I$eCc#���,`���Ғb�x��鷏Ι!Ձ鎆�m��8�})YK`���׏�H�X8�� #s��W=��]�&A�r�I�v���ӻw��	( �SNYs@a�@3��^��4�98^��)��y�
��^��L*��8�/�H�g<R/ɓ�Ӧi7����~� �6[���)� w8���S) Q�OV�@�PW���Jqo���c�����$Խ01�ޡ�a�p٫�y
���@�nI�E/�1���-lѳǓ�}j��,�Ny4�
��>�!��'�J�3��Q6U�̸'<�<�"e��5;N21֚��rH��G�np3���.H������ �@�)[=9�R�b?N��8#9�r� ��yۃ�4|��i�L7,[9�);�����	�ʚ i*[��g�t��?��}iJ�� �6��g8#�֝�NN��E0���8��S���<�4�q�{P����Q���׊8�9���;&���zR������Ӟ�1ޝ�N3�@�{~4b��"��Z 1��݁�2��Pm��:�R�݃�j��'�7̣ڀ#*P�cA�s�=6���np=)U�y�) £�~�zw�hݵx �_��<SX����)?�rE2I�@R��ҝ�.៥&B�CH���1֓���)�T���4�z�� O t�+���=���e���Ґ������*�ڕr,/Ҁ"�˒y�]�eY�נ��s��m���[_ܩ�B��I�Ō�T"��}:׹|f;~ő�`q^�
x�G���7�x� ����� �<�(z�r?¾�-��3ZG��7�䍱ӥlY�CR�;R&f�@{�� ���7�C(-�z�{?�������$UƥGA��ν���dyp�uv|e�xR�Kb���A�aֽ��%��H��bq��� ^��#�zi�u�P����Xq��y'�;��ȱդ*F>���hu}�&�TY��������јs�
s�����&+ʙ�#�j�����D�Y��k�Eo�N�|�h8$1��f�2��ϡ��FP�-��##>���˶���fq��c�y����_����+:N�ë�ns���_B|�> �ʷ$�ޜW��bσ���{��#��	<I	�R_β�uCc��OH �P?A]ČU�l���A� �J�1���w�ke����擎:��J��㯯j�a��p�Н�1�WP�]Go�����7���-�����u��n=2N+�Ե(�Ī�Xzo�o�	ݟ�+�m���ca��q�WGS֙�Ku8�,daL��>1x��l�_���ӆ�tג�	�����Jm���9"���=&�km�h��
�5�U���h�i;��V�������]\���Kk��*�'3g&���:־����l�?�$�ڀ��d���A�G���E,QO�k���<I������]�ȡk&)��zW��n�eU�w`n��_�|'x�G��!����_L��.'o5��lB>>lξ��� Ħ3��(	t5J徕��C����8�,�ƨkr�vlO��"O=�5�H�G+���1ZZ���wWy��KRb��48��5@s�

{hvm�c�?J�?�%���RpzW�[��j <��6����1_|PLX�:�ԣE����V�G��¾,���K`�tg��EzƉ�	��6���u����i���;�a��^�{=�����>]��r��b�-ϞgMn��#��:�ʞ���V���خ4g
�8�g����ukO5�ɴ�v�CT?�u��+�q�L�[���ٷD[}��+0�����.�m�"���@���?|&�^�ev�Q\w�_\x�^�)(҇���^w6>ڲiq7v
O�+�Xƹ��~��F�Y�j��Nk��6���?�?ʽj#�ג|n;4;�zm?ʹ��T~#�[�c'������|1����G�.+���p�. `B�<
�<9}5��<y������T�&u~$�\6���2zמOgr^v��|Y6�=�H��_���滑��7�������)7C�}K��Oe��b�Q��ߑ:��s_U|)��V�#o��sx3׵K����+p ���g��}fmQ�\��d1����V�~��q���W�:���#(+�p��NO#���rEٟ���+k�c���2d~\~5���3�-~뺼�W���J�y�#>��?�.�]?º��$D=9�� �Z��ۃƒ��8�e�w��x`�H���GK��� ��|�X,�@9<`� \
�	���,�(��9\sۊ���!x�N���I��ҿg?f��|Q�kW���X��\��֪���6����~3iw�g@��X������u�J��$�s_�� �/�`��/��b8�L|����_�4����"��V*=85�e�NJQ�s��n�W�Z���t��|n�r61ۥz֟��P��kP�_��)$b�.F@�U�@�)M�{z��4��s֔0ϥE��S���J szL8�O_Κs�j n�~T�4��<�Пz��>�0�}i좐��@�zjua�ޫ�ԂM��>r��+�]�hW����<+�ǥ^)h�{�l�=�:�Eݢ�@
v�{f�o|d�<;B�� q�zc5�E�-ZG�xO�?�,5K{�.(�Vw��F{�Q����o;J� ;�2�ϖ
W �5�'�%�y,��206��~b��^׮�M�M�]�,���T#��☴���(�+����My��H�xR�#6���OQ�V��/�F�+`z�n�����^X؀+#V����i�7z��%��p�I=iY���Y�z�y�59\�}�&��Ձ,r=������!�Iթ+4�;܁�k�����z�@��� zz�N,d��5#N)۔2�6���1,��2:�i�\"|������e�T)�����:HA��� Z�A���({�����랴�5Xs�_� �޹�|᳸�'�Ξ���=8<P�j�_�8��5/�cR�x��Q,Nx�Ҝ́I��4����n���ӯJ�#��AQ����i�aϨ?�oJ�����v� �-�����z��[��>�ğ�Xn��Ѥ�A%GO_ƶb����,��On?CHun�92��7'���m���5��\�9��5�k�y��r��x�d�ky��v�rv��� >���]"������^Q!�v�8�}$~��FY ��pW ��5�[o�mv�B�{,i�g�J��o����1���6?��'v8�n~�h�Ƈ�ʩ�Or�u�֬j;�f�q�D���G�׈�J��9;�#��C�Z]��f�������wG鷈>$i걄��?/�1��x�OH��_���l�^����&���M�5�� � Z��;֮!�&�]���<~F��пim�\���%ٶ���"�J�f�ܪ�?+��.b��[iѾ�z��~��ڕĳ\yҹ�f�Ϟ��%��s�6U�'�����63r���� �WQ�v����6&���/�v���;�x��x��������ߘ}=j� ��}jf�*F�U�(�ue/�#(�zt�|�,�pH �n���Y�s�}�	�r�8���#���r:SaPː6�h@��9�8���׭P�t&���~t�>��_�s������I҅o�ۿ4 �w�3Fߗ����I�^Y�8�
(x8�ьc�qQ��A'�;<P�g���}}���Kʟ^h��y��QJT�����>��($�� Fp}iy����}i�0:z����<R�s��T��~�}�
�O\R7m����v}}�S6�$�s�;h+� ]ŗ���M�?Zq]�{� :k�.�;PH�P����r}qI���I��#I~�+���( �3��G _4)h#�1�d醤� ���� � 3n�w9���g�4�����NeH�=� [��NzPv�����r>��r`~��sc#�}=���7 �{�$?ÊC�W�00��g��K��(9��9���<q�U�g��>����I��>� C �s�P�!Y�m܏����a�`zf�	8�=;� ��fV����C�?� X7�N]~v���TNr����)���<�;z��f�h�@RUq�O�4�,�*�	����H�	��Õ��dc�NԿt�)P������i�;N:��o4��riy4 �bzt���+`. �- 7�8�Rzs�z E�?��rz=��� �F޸횈�����piCu��׮z9nOOj_,����n!�2*?�R�1E~��`�;�4`{
 #�җh���� {ڕx<i6�ڕ� �Q�`B��SF3�(�׽&�3�\�����'$u��
�#�b����R*� g�cd�9��R��3�4ݻ����v�I�>��h��� �4�n�8&��[�l�r09ϵ ~n���ɴrG�&��-�⍤�~�&����)&a���� %�q�����Á�1� ���[��k���Ŭ�0;W$W����;�@������6� ��8�\�ǃ^��zE_'�ea�����^��x�!�i��=��W��W`�I��.Р�Q�����˞���O�3��/|���6N	�Xc�ƽK��%��62�۽�*�CᏏ"4��J�󯦼�Gg>�>�%�ϏQ��]����V���~��� ��HT���S��π��z��>����'���J���~R�ջzW�-�oW~2���������'�t�q��V�|���~l��Ԯ��ʒ��<9��~�x�?♹n`�L)ο2�E_jq�}˧U�=����������ĆE8l�߾kf+����$!U���������۸��s�#��\��7<3��>a��#����m��2+�c��1�����#�쐩9l�����\����|]���� �-s�8�+�c�{��c��ғ���zQ�)�M��������wJ��3,d����.4���񞆢Ӽ:�w�C+6{S5q��F�v��ڕ����X��3��0���z�X+c�j��]�=Xd7��G�|j��^���B�����V����$ k�?iI�i�FFY��x=σ��5���Ιi]��k6�����s���׻xz)a��\��j��~��B�"��Ԋ��A�F�)-O$���M���2Fx�CG��úl�a�$�>���3�s�5�?4�n]��ԍ͌c��>�w9
پ��u��|�ξ��mŞ�`���;�W�q��.&\�#�z\�l�ا�[����0��q�sҭc�Q+BwzT����(-�Y��5Vp�ƍ9+��K��>Fj|1n��W�<��F���&��A�p.�X;ȯD����gmyֳ�I|�*��� �(�`�gMk���a-�`1���MKXU�e��$�wZlN���p;WC����:΄��H��K�YdZE]�+����l\��@�����A�[~cM��ּ�Y���4�E�H�<�����T};Jc%�g���5�~&���\�\�\�[8stE����H�����w��:�m��v� �_=���:_�<��Y�n�s^������Cc�3)�>cB��r�c�����6{T���ud�t�p�ȭ	~\��f���y�����a�U�p}�Ƽ��km�/���
�Cs�7�u�:��w�q�Y?⷗[�g+��7t�k����5K��w�^��8���)�j�?	rճ�?h�;�r��,j��=����E�:�ϖ9s]W�5�zk�>����diI#������[+��G6��σ7��P&�( c5�v{�H�Ny9�x�G����"�{�ZP���[��)�)��_x��l�">��8�%���=��W�Q���G㶾���	�xǋr�d��oVUʓ����ˎ�Z�˾0����i?!�Jp	]��׎��~%���&�f�~�����v���J��c��Λ$m��:�~'|I���;�G�rO�K]���o�s,z��'�}��W�n����6AqfØ�<���?�_�5������+�J���F���YUKcH�S�~'��ڿ��	�V1nfR�'��?Z�[����;�33u�^�9F�y���d�x�v3����;�[JВ�$lr�������R�i�H9�g���#F3��Cwe'���R�fPUh�����ϥY�@���搄�G4��qSI	a�ޣ^�} ;���H�n�׮{S_�Ȧ��� �l6���hPH�F\3@�M0�^�o9��Q�q��Pϭ+R`��:���ʺ�/\~F�^L}�U2y�j�!c��¼ռ	�Im%�\ c�c��W��p��X�]Y~_gh� �u�
�����ʃ,ǧN�����Ͱ�+vt#�+��σu-|702�:����(��O�����O[[;��Nq��\����cGUSW�C��
�<ct���߳��� K@��E0p_�m�FF�F	�+�~'i����Z��C��$�F9��G���Ws���R�Q�<��}&���*d�t5��	,�&D#��q]��Ժ���X?<n �z��*4�t���]��jr��3E��PB�d�9����>hW�k��n,l�A�]��U}�w'-��M:Fz g�f���ku��L`�� ��cJ�uu�]�3c��2s�O������>1h���i<�Uu\�z�_@|p��t߆��t^+��)�;MMQ��bWʜ&1ם���ڼF�nl5�*h�kpd�h�3�q_L~ӟ��Y�;��(-��+��擝�;z�1��1��R������ӵ��A�ߞ�}�գ�|��8���\���L�s p�I��
��|]�I#�B�璸�=��[\��U���Ò�C/�qYrZ�r�#�ɯ\O�uc"9�qR�N{���q�:U�W%�fIj��������n��N}j�i��O_j���8$�߶Oj�*Iy��֕�Ѝ��*`ݖ�x��UY���ơg�V$��u����U�J�e�TfS���8��-���s�N1��]�6nʐ0+���� *�q���M;C1,�����d[��ޙ�j�ڕ�
03�U��i0e,��*pZ��|��p���z�jJ�vV�����FC�'��� �2-&�[�9U��n�P���x鎄�2!e%Aӷ�2�`��L�S.��H6%�1������̂M��*O���_Z�!�@�q�kB6Y�:��@� >��h�P�n���#^1�N:����GK�����PRx��]Ή�-�=�w��ָF��w'��lgӚ�,n�ceL� �*z;��|���ï�s���<0�\���9S��ۏ� _�X�IUN��Ð�?w�>�=���>�Ò0qO�+�v� �z�$ M(���Z R}�I�Q��м�GJ P� �ZA��~��7d����� v��z��J{��Fӷ=� ������q�Ͻ- .}�����ۭ%&~`;t�� s���9X�x���A�K�7 �l`��)��Ѵ���zӟ�r3�曕�Ҁ�a�70)<t9����9���4dzq��ӷJOA�PHq���P3�Z]ø8<SyNG� �N8����K�r�{sM;N�z��R���J0$�b��ozRŤ'<d9����� Z�X���.T�}{f�*8稦I��=ǧ�;���@�y��P���v���zS�ᾔ����!�~� n`�i�m�gژ�n=�� ֧�� }��Veت�q�S6��JDb˓�}i�z��zP/ldsS�7�b��rj�l/�E`d���'�`_�5������s�wϥU��{�m`@�ߎ���?
AR}(�N3M�;?��P���sF(��q�sK�zRn�>��4�SA�8�(,7c��`3o�ךwӚ_\s�@��<��4g�p}�(�n�� �#q������S��N$`sH�v� �X�^9�	����q@ x����4�M�9�5'=� �R =�4n�qK�4 �s�Ҋo�;�h�׷jk�S���ޚޔ�5W�ܓL���9$�jI$ؤ
��ks��,D|��Q�x �ޤP�z��|g�8����#��p��}����р�$��P ���)$�r�������Hƥ��s�R\�r���<�f�i�x��h0ߝt���T� �¹��T����à4ynG_sM���?.�C#���p����^r�=y�1�f�_���A����� �J��:�;���@@�*q���6-P�sW��d��>L-<P�r��8#�f�C<7�M?�D#r�:�*��z��O�"�����+���ޫ�_�G#}��w��c�WT(ᬏ�i�Yu� [�$ޱ�mA��X�7͝�H� ��^���~�\\5��&s��u:o�;M"�z"�(�>�_�J4��&��~3�D#�n&-�.Np:t?�~x��%�59"<Ip��7� J�/���\��X[K��+`���b�d���q�b����J��|��?f�Ig�,Lx �}�	�k?/Ҷ����� ����-�U+�-�_C����hs�¾v��b@�;�П��փ��t��:�t�?J��R�����`��O�m�Ga3�»��7=+�l�~�v���R+n�ѻߚo�9ʀz�@ǅ�*���L$8�U��@$�%��cf���@u)$��;��9;������ֶ�7b���r���I�j1�������S\7���������	�r� �M+���D�h�W�W
�^�ą����mށox��5�'#8�I��4 �����墀)7g��r�4���$Vt�Y�x~�{�#�j���?ʟ��`�c@��"��$j�SY�=�J۠�h�&���j��0�������v��%�#��Ў:�\[{�����/��a�\ן�β�Z���9�l�>�VD�GU�!�[C�&���lua�y�ݻCx�b���":�+�Vʹ!=� ʹ՚��8X��1W�?M8 |�޳��=�J���k���K(�FN�XL3�񿍺���ʀ�f��<����&�p�<�qL�y��� �Q�]_] ���#���+����_�;P	d���������N9rx� � ��� �!0�I��1�P����%�ro���g�xf�G@d+���3�w�W�:�sڮ�BNG�v� �Mo�x~��	��\� ƭz?k��w����4�M��{7�a�s�G�+�&��^_�GGkM˴��W�J�y�}�ń���:M����W��޼��c������U�[b�����+�Z�c���[�ڥ����G������W������5�xK��jI�8-��Q�{���~�d��EU=1ڼv����g�N+�|Y��W�fH#�+�ﴃgpЌ��MJ����X�[{f��׃�k߼��'B0k�t5v��Q��dt��|�F���;�s��4>��Y�(�E���d[�V�����+�>9x&��Z�r�t����JഝZ�A�}���[a�uv�]	�H���*їf�ym���n-n��v���x���M.�H���x��$�WZ{D������L7�]�'ҵS�Z����;�i p�w��k[8�@:~_L�����)��5�#m�p�+'.a�E%��`��$�+?�i�re�|~�V;zƦ�Tm�x�ӊUm���+|� ��)����(�/\`t��R;�ʫ����=[�yƐ1͹�5�@?Rj�Qޜz�����P�n�G�H�01MV=��3g�qCd��=){(�8=G� 4��1�"��4�0-�oj�9=;��F;S�1���,��=������S�m~�6�p:��u��"����h~y�C2��c�t��q)�5�¶ 
w�aֻ�Oh�=���\���"���Z.�����> ������D\�De�����	�K�Pi0�w�G�����FA?Z��#|F�A�mt��B�������`w<{q^]�o�M�[]2�!��`��� ��D�A�͟ƻ��ܾ����4	:���,8�=���\�(М��.��9ϵP��>ta�9��kY��(�I!<��ֱ�Iܮgk!�;w9�#}�cN��ǻx�wXx��t��=�Y����p�+ɫ��G"�S�~uF�1R ���SM��@l���Zض�+ ���V��>&��&��Y:~���YE��+fKԺ�88�Y��)��� �R���׼N���G�� 	9�w��g�dړ[EvXC��ι{�V���#�&����Nzҗ"e9;X�����`Ͱ&A>�޽��}���Uk�J(䷄A�?N��x��n	`�ǰ��+��ll�;FÍ��>ب�>m���G�^<�|'g�멦ڬ�#}���du���n�]u�`��zqZ�x�Ph¼�\.���5�op�3`\�q��*)��&N�;8;� s��t�e!I9���%��a��������uY��+r=b���ddd�p~��5��"�\�z/_�t~,�������+9e��݃�~FG�V#K�q��:���!�ӥk_F�#��;�=z�U��\�~�B�Ӟ��3~�����¥�1d�tE�#����q��V��B�}�W�.���w�E}2,e��!���t ӡ��|]��\$zf�z��g$s�=sJn�7�U�r���[�Ycu�WC���C#���}0N{g�W��_�e����d�?���|9�վ��@��H���RX`�g�4��.�b���|?�/�6>Waߥ{O�� g� ��$��̋�0Tך��]�|?׾�_X_ĺ�p;[G�lc0������'�_�MW�� M:�ǔ�wI���q���J6��/���\?<eo5���ڃ8U<lq���ɬ��Z��{�+y�f����:W�~ܚ�~2�Y�ꅷ<J�������%u���k��`��FB�WL%x;����t?�Q���1E��n��'����1|+���Xq9��a���WQ���n��8h���2�����YGw���a�/ `��e)s$��V<�Voj̮�[�q\°�����\%���/��o�q⸙�ݸ����j���b��'��~�7@W��jp>b�kB@~�[���<S��v2Fz���~�E(�}����=){u����^�4�=�43�<�6��N�����H����� �$��) =	�Jr�ON����� ��/?�����Ґ���-���%/z������(8-��go���8#��$V���Z �2��E!9�'�LUNq�2�:Em�R��FF@��0��� zR��S�;OˏAHC9$��}��{c֏@�ڎH���B:��i��$mȤ,p}3�+}�}h F±��
J�H�=zRm'�?�"3n�H�h7NI��4n���7͆���J[,GA�ޘ
Üy���y8���2�׭=���i#���@Ŏz��Ne݀9���GLS���{R�m�����8�҄���=����W'��R����1T�-���G\6q@9X��vrN8�F��s��ڜ�Uq�ۚ[���;FSB�>���Dm������;A^G�Lb.{��G8�ځ֤b�I�zP��h�ƪ�l��ҕ�8?ʥ�B̋���*歧-�����2!v����ñ��'��J�'����P���#��
�X��zk}�ANYyA4y���LB����& ���{u�e;��@E!]����"�� :(p:���u⌍�=i�N1�4��Q��:08� ��V=���7����� �
�:��*���֓���ڭ���4�@S�څ��� /��!9��� c�Q���@���`�����;Ҳ���0�a���㻒G<�i�S���O;~ldm�}�W=s�@4�\x�
On��e?6zH́�� �s�x�*����߿����,0)�z�����ÿ�lÜ;R�9���2RCg���0��t�eB&5̶0+���#'��4Й�xSX:/�#�T>?�� �� �M68ь�F}+� ���L�}5�Köw�f������sh�GV{D~<֯�2ZX��6�=�p��-q�ۓit�;�8ee��_ex7��r�lq$0@��L� ��G�~j��Zm��}B�IlZ���*r7��Ǳ�3Q�\j)_C��i�CT}����6����4x���m�hc��μ;�φ�37̪z��_|%���w�Җ�J*���zP␝KGc�S���j���&���� �8�|,\z�U�� �sR�t�mC��[�B9sq,c��������u�G_��顕MRe=�g�x"�HA��w ּ� @�n���'#��g�љ�gûQ�~z�����E��ϿOҾ{���'�z�ຆ�=�S�W%k�d6?J���K�?�"��rsҸo�_�rFp�ʻ�������3��9@Q�g�4�v��y��Q�\׊���G���Ӗ����'�d�BU������i�³���M*�s��;�E����=�ۙṾK�ٵ򤜂+_O���$*��zM��;$T\���t#5KG,4�c�굜�?	C�s�p:�C0P>n:
��u���X����5�6�w0��fϯ�ې��`�N�K���^w7�mkQ��l�AJ�Ϫ����n\�ƴ!�I�A�������ַk�ȭ�J�|]R$3��}M �֧��w����Y�.��
����h����-�bx��s����<���Bm=�q�&��5��R���	�Z�URE�O5����t���7���w�Ԟkx�X� �Hܠh�@n�v���}І-���t��B��k\�)T��;�$��uD�bw��ֻ{[�:�3^kc��ou�I�O�z6�-����+�ed��x�'�w�ε�0�#�1*�#�ƞ��E$_z�����_<?��I�)��;㾛sy�]&Ӎ��W�^I��� 1
yĿ�jQKt��u^��m��G�:��k�TY>O�7�⽧���{�cUK��i ��s�:��@�!,��G��,--�c�_�jP��������j�N*�X����p*��w���^U�C���?�z��y_�O���x�z��͏�6�s����=����F����~5��FP���x˜~���wJMWVH�����5�*[��|a���J*��1���^�-��&�'5�"�-�6�� N+��-5m�U8@r�ҕ��4+�2r%���< ��lO<k��Q��[�����H��:*$mݼḵ�Q"�m�/'=����f�����L������}/����Jy��/��� :�~/~��n��Kk��I.�(۾\b>1�Es(��gr}2�����e�yR2�>����m�� ��|���z��P����������O�_Ǔ�Z������0Z��l9�y�|M�`7_�`�B�ՋX6;�z���^4���7+u��������H�Y�<�����9�A?ʤi��p+�{�^*��(�k!�����I�T�mˑ�U����~��*�?�3��)���p�{�*����*7 ���NfVQ��*@��l ��P�1�T�S��;�¯B˴�y��J��b���5egڤ�`����i<q�Rϕ� �qL�
���Z��0�t��q�9� s���z��D���,ۻS�$1ɖ�)���㊴6��1����c����+:�ᝰ�T{U�Ղ�@�)_+�'�v^����5>�� #
_@q��rr8�.k� �Fd$�7<�m�i<'�u) i!b�����8�:/FS_��XܬJd=���k�~&k� �O`�c۴g��� �k����t�#yc�f*y �����|��8%�q��<��w���v8t<�S�s������f�3Y��[�
NZ�լ͵�+�s��5F�8�{O��B��?C�+����*3�zΟ��������0ߕ+���E���GS�~^������$��B�������'���4w����^�� :��"���ճX��v��x8Sc��\���ր:k����rG�|�ӵS��x��s�ҩ��U�Id\�F�����O����U��#Ҟ�F8��.�� #��|z���M��y$����������O��R@G遚�=�&�*ۺ*]���<dw��otr>�&���B@n�s�0+��9�MV�f�o~����c?�ԑ���d�^�i�:�و^3ӽA��\�F$Pԟ�B��fe�Eg�I��<:>Q��������[X�I���k����Rzջ��L��?�Ӡ�}je~�"�Ǉ���񴐩���G5��x�N���o|��H�̅�q��>� Z�&���bT��U�|2/��cx�0U�	'g�d�ʽ�%Ҽ2�xF�nݐ[��Q_@|�O�k�PA}>� t��z�>�6�u82G ��a��o�5���g��R������R.��;�S|���ɢ�d��ak���<.�Oj��~�����\�Y�`PW�;s���W�~�;��],�I�a�z��������x¾���;rYC1f�N��(����5un~W�֖�h_��"D*[PB�T9�f�K�]��o��*�r�.B� m��c�~�������=s�Y�[��C����f�>�.ڂL�[;�9��y�8�V���F2�����ϫ� �2+�-�H�J�����ݽP��?�sT��xDR���r�8�O�fE��2�˸)��ZۣD�0��&h���3�r��1r�����w|�ɮn�>f>�/ִ��77'�A�GjR$�4��ʑ��D�����~�ǭ!*��98�sߧ�( l�.GzV�H�?ZL��n�%���	 ⥾��YSg��5rǌC��J(�QH;Nzs���������q��s@����*���Ѵ0�=�.��Z �݊�QԜ�a�@s����j�Aݜ{ӛ,� 2���k=�y$-���N���<�'OZw$��~i�\�.G�jr����zu�8<q�)���l)�{TΣ��
ac���� : �ha��s۽1P3e�<`b��F0�P2=����ƂH{FsJ�� �z�5,�����H�zP�#�~m���L���?�4�=��5#õs���銟�9�}1@�>l�ހ��G��jA�rUFsO����}��L|s���xܥO_QRE�,�ۊO%��\5  m���q��ݦLps��J�o��ҵ���%��Z%!W ��u�m�~S��Dm���͎hPv��j���sҤ����q����k��8����rF1��� �����;����NԁKq�z�ڎ�)�/p(=�CN�T�z� �<P��hy�h�gq�����H� q�S����4y8�0q��j����9'�՛��h����(#�@�n����s���E��Z?1FF;���x�)rc*A�Fpy4���F3�N��r9����?]�@ǯZv \�P+!���zU��gҝ#s��r������Iր
LJZ( ��4Zn���ZQ�ϊJ_�O~M ��=>��I������� 5	�� ��#}�3�J�6Q�F	㞵$*�̭���@�c"�a�B�x��O�6�|���S��rI���L
�0�=*����EY�V����叞O�&"=Î�09��j)�{�z�R7��J�w8��OZBq~=i��~~������Ҙ:���z����e�i��S��^}h�Py�����֜�zdd� ��I���4���w\�[�9>ϵ\eXg8�\�\���;1��w(��^��a���J�<��_ڏ*&�q�v���7��y���u�ǌ`�q��Ua����7߶g�&�^��ᭃ!M�E��^yys��Rj7r�-܎]ݏS�� Z"�]�1�qR8O,�@�8S֒��]�v���s�Q��y�+����<Kie���kud�$��^	h͎2{s�����
��Ni8&W;�c�^.ռs�ɪj�msx�>cϦj!q��2q��x��/�0�)y╰Ct`r2��ZV"����r�����;�0��� 8ުN���� ��`�{L�7�E}�O��5�'��t�F�	=+�/��V��ֱ�uCc���Cg��*�NO�Ҹ?���.M�?.+�<��Ͻt#bs�җ܏aNc�i�t�#=�0�v:W;� 6���'���\ǋ1�!��<���G5嬍")S/}���,���^G$������sK��|��\��.����c4r��Ȼz�c���H�,H�W�a1�Ƥ�Տ�sڂH�$��H{v���/x�����g;B��{W�.�:\�q_)���ox�e/7N�Z
�ט����~.�7��^V9 ��21�}��=���ڪ<jX/<w�/�zZV�������cԴ���:	rrg��-Ӯ�(��pW���|<�ó��9,:��j�y�'��x�A�T�$;K�*{q@��]��O�Ǔ˶�� x�m}	k2\[�)�"�A����� ��)>6�k�_\��I���	�Ir��gi�YZ���ف<Z��|�k��C`��
<����P��(`ޙ�$q]� ��T�[�h5���_M'�y$���"�b�<��4�Go*�p�(�}�^o�.�2c��z%�Ŵ�����ϥy��k8�&f �\�ށ���4P͖�y�5�Z>��4h��q�^]�٤�El���^��}�1�ْ��S�հ���e����m\�okQ~���@�}��[��O˞�u�N�ǒ�_��-��ed�K�8y���I�_\LҼ�"�8"���_��2�.5;�û9U2s�ի�o���4�>�n=�KF�J/��}w����e��r;v��I�v�����|�sS��{i�xn'��?
�>,xT�7Z���]�?;h�Eu)Y�}���ɫY�S�#�T�V5�5�5=�F'�E<���5��7͊�'����30�Ⱥ=>S^�k��2� ����cWb�����3X���^wc,����X����fN�tO�k��Ė�"Σi=�(�%>����[ɬB9m�zן�^I4�[�}+��R�]���"���cڼZ�hd�ʨ�Eà�[� d+��5�
u��R�N����x�6�4�g���_��{k RV�{���ձ��j�?��Ҿ1��p�������}��d_"�>N?*���iǋ8�� �YCr��cxT�D��Ⱞ셔�ea�G�}�����������;#xd��Sb����񨛱����_���5d��s�NzW�@��@�~U���ӪD��`��9�OҾ���|��x��
��Y�� t�z����8I�������;q��.���
g��}���Z>�o}aB���� �����n��^�f�	� ���k�>�WM]M��\.��*I��V���2@#����+��;�������[��q���h��zNU,���[~��x�z��� /�a�����@�[w�:9v��Lz�m�j^J㯽I)�r:u4�� z���f��'�zԋ��q�Ҥe�x�RIɫ�@��<�UVm�x�ր�i�>81�~(i�x�}���sMb���98��Qܹv�ߨ����ペ�f��P2���b�9�����l�;�"�W����n��ֽ�P������/��*�g������:x�*x�bPo����,q�l
�uV�W�k��.�ws�3ޣ9e�:�B�1�2� �?��Y����c�.�|��'<�z�d���1&�К�7`�d��J��N�gޥ���b�ZƄ�\���x/�2��g��N�vğ9��V�L�Fc�������V�����|�<�*��2n'��?�X��i��1�^� �Q��\�z��$FU���w�����ҕ�h.\�MX�9�`"� ��jݲ�0��=G�UJ��8
9�#4�R��@Kq��8�ɩ ��hdu����I̖���I�ƻآ����=��֫���v����[ǝ������ت\���<�)�j;�<m�=��wV�Gl�rx�\���i�A� ҉�>���3q
�'���5�g}�;�N�N�5�NN;ԗ�l�RX�l#��omn%��bf8c�z�Q��"��*rx����'����,1<gzU���jF{��]J�m幝\�n`�c����-5X#�-� *'��W�.�ug2�h�NO'��R7�o�&�D��L�O��H���V+#��P�#�"D
99m���@�恦\0qF��w��~enjJr������ޙr��Z�`� ���9���u.-�D�r������G,w��1� ���Y~"�ܷ��Ex��t*0�����8�i���/ˎ��#ۚ,�"�;;Gy#J��׷z�ٳU$��?j�4:��e��`TQ��μúM���ݮ�L�*�N���1�c�#�u��Z���Ist嬏����滯�F�=���NA*@����uq�)��1���Օ�B;Ǹ��F:����l�(��6;�zֱ�Ņ�`�X�ձ���������x�Ve�򜎼S�cH��#1.�Q\���pMt���VېWo$���
�x��&0�y=�@�ȣ=���;
��SKA��v>�i���)�Z@6)��4`����Rs�J b�������������@��:�y��!e��4u�~h� "�;u=y�AQ����E!�돥 '�Oj^q�	Z#���Қ`86��Jac����F�('�Q�H�� �;��4[%�g�F�W�)~`� {R }�F?�j7���ۊC�O�W��L���lzz���e�?_JF����sϷ4�H�<w��SU����HD�(���3�#�:Rnp�r��c���뷀c�Ni_����s�L	$l/�3ǧ�C�ߝ7��9z��Ԁt�՗��ȭ��4˗�`�x��dsX����7 h�ᤍ�����
�,/B0?*�G>X�ክ�C����p� >Q"���s�lj^&���cҔ�۬�kc���~�k�[��4��FKc����p�Ђ:��?�,���.O~�m�c�����ʫ����H��J���\��p)�]���֐(V���c��z��Ps�� ����sMR1K�LQ�Ɓ�$�z�ԁ�H�QK�v⚣h=���3���pOa֐.,✹�B��ֆ[�d�)�J��{���ǯ�.x+��Q� �S�O^s@�1W�l��1Ry�2�ch�Q�s��k͞	���`˹�Q�S[����n�y��w�
�q���q֓hی����+�FG4�U�Ϩ�Z	�RR�z��(�aKHX���I�E8c��o�@�F>a����B㩣�A��	��1��5'��e*T���UN��=i����
b$� '<��V�r20{
�e;Gl���wA�pL@���n3�cr��+a�<���q���5 '�	�):���w$�_��0:���~\P���1I��NV���� ��F=�$�a��v�/�ӧn)�8�@g�t��,v$��\�u�T`�H�,���q֨F�:c�j��Yw^RJ�s�*�Sm_o��Z{u!6�Q�N�{;3sܞ~�B��#���M�S�>��(ef a[��1�5dd'q���Y��y�r��1�Ӛ@0��	��̑�����j�����r ��M�O�嵩E�ɿ'J�E\����'�:��+7���zb�.�y��v���?X������;c]�U�=:W�>6�9�o)WfN=(��1�1�i%��{��kn�5�=�x*��� c��5�� �#��݀���?:��G]=���� ��K��ֻÞ�+��F��'$�z��px�[-�F�g�*���m��%G�>�y��Un��x�vY�`޻:޺��8�ް<D����#=���~�5	��U�EC�<V͎�Vf�b� �M���e�>ՒV�I�I���5��Y}��@�K��i�՛�횸���=*;P�f�Nx��6Ǹ�����;^���P;W�iJ�_i1qӷ5�{w.�Z���+�9�@]�l�K4��F?Jc^D����f��ş��� 32��5����gf�36���B�Y�^�T���It�yi"�G�5���C[\Ϊ&o�^���Vڣ 3�pz�K�DZ���7ZK�F�Ê�_����(���V�o-��(Vn�>�h�;q��x�5��[:���d��;x�*��ʰp@�#���SNf��޵kG�b�.�!L�a�q�z�1�˨�/� (���߂�Ed���A]I�6���W��=.�c#m��+�W&��8�����K��������#�Z��@p�kм+*[��,1��1�h�*���ڷ�?Y�T'4���/�(��?�З���v��^��H�^y�kãV��dL�/\{b�1�J�~ΓD��[ƥ��g�?O֬~�cM�d8@� �Њ��G�'��� *���� l�.4I�.��O�O���yr� ��|3 ��X�}N��kㆨ��}�||��5��F���"oݶ���[�O�u/��}{�!Z��r�$���� ��,�x��
�ʽBo�j���u�4ԏN �r6_�#&��"�+�ˏ�{��O�S���ߌ˷G�� t� *¦���_���܌���4}6}J�R��۫���1�]�݈��X�M�#7Bn�޳���7|A��V�M�M�����1��e����Ӛ����:�g��B�v��u�b-CS��d�J�r���eA'Px���~��GlϜ+�YW�T��_E|-��iO��(��A�}3�F��~_9_�_|W�v�u㴊�7b���'����I�V��aZu�rA[��g���w�_�F���ݬ���8��5����������[�è�ђ�3g���/���_�w��H�j�g���D��t�
��8 J��֬5��6�l�W���8����R>`�Gc)�	b̬� {>���7x���M2.��#�|�������,��?2�u�ǂ|:��M�4a��wg�ִ��d��{� �>/h^�}�[��I����W�ƭm���j%v��wO��W�4�^�JH��͑��@��_/|M�h���j�{�ec���nb�2;��e��̼�1^��h�c!w7eZ���	ۀ�+I�n$l�Ll  �+Ed;@-�ֲX3ciɫ;���ֳ(���y�iʻr �FN���aTn�&m��*�p:���8���;T�"�8B1�괨a�}G�9�h$g'�M*�]ǚ`E$x_�H?J�1�5mX/������#���
�g�Nz�Lh��l�@8��n�����&ە�ހ>]�%+i!�OʼJH�;�VN$��G��{e��f o�Y����^;.�}%�1����λ�q��VU팑�V�t��F
����}j���u	�EhA<+�#�x+Ð���9����*۱�������;G����T��g�� X�9����k���2M A��n�a�D�`��i}`#��?��F8��s(��y*���*ũ�����w�2rJ���Y�s#�V�����Ү��?)F�A��l�F_w Ӯ�������*e���۴��M0)��Kv�
c3l$g��`���O�J��̤��?
`*��"�v�Xt��3�����~���KF�g�as�{�׬�=�^�u�jww/�-�ٰs�� YJ��Eƙ��z�a�I� e�if�����#'w����E4n��������T��喯
G~d���i�	�$v���s��R}�� �.OR;ּv.�Wvͽs�Q�Y�f)�ld�ϥ]�Eў����ңef^���M$��y�t��5W{
�c��c>\�ZvZ�kqo0TmW�aT�v�2�UWvV���@[�t�/1������xe'��]&�p�
c�o��5�}f��1Q��LPЌ��pZ�&��9���z����T٨|�Wi#�P2v�-! ���N'�X����~��fl~�zU���U�2�Gz �h1����
v�n���5�˵�t=UP�~��V���%�E�ҋ��6	���z������.��(�C���y弄H%'(2k�<3�Z��t��T��E�FW�:�[\��<��u-ԅ�,-�[�OJђ�/.��&�p9�)������Y��6X����ӟJ���k�y�܂	��:�.�z�>T�^r�ǹ�f�Q�z�޻�[GY��m%��v���kֵ��I�����[�g�+��p9���A3�6���}�R� �8��H�$��=q֛��$94�x�C��Ca�'��QҕW���S˜�w�6�;
9�{���L����:�R��=�BpNz{R5b�����G9��x��ˎ}� �B�n�:
��M+ ˎi���E.:����\�H��1K�#�;�@	��R.��V�\�?�Q���0ޤ })pY~n����q�JI$�@�^s@��Q
��-�b��V�F��.��c��#F�gސ�����F�Ҕ��>_��Al�|�
�ys�(�Lnhב�{�YJ��8�4�����W+!�>��i���]�h� �N?t1��_�	������?Z<|�·P˸z��$|�(@� b�˰8�����8��9�S� Lc�ґ�F3J����J��ۭ H�� .�sґY�eRW�ސu=���U�G�ך �q�����~nFM'�$צ9�0A_riN���G9ϸ����0K�`�5O8�H��#Ҙ��;��e-���4n<R���H\���R.���4��� Jz�ˎ��nN޹46U���?Z����ǻ���(.�U�H �{w�F����H���`{���<g���4w=��4������N-�FiT��v�`1G�A�_jC�I���L��?�G�p9��f+���L��FO�֞ܨ��&ߕp9�<pi �^=}�����e܀�~Z����~f�1�b�^�h 8<Q�-'_�@i~���=)iY�6q@r��ҐbNO�K��Q����!��z�S6����O��pF�\��� H@��ܖ<:��n8@��p�xp;ԏ�_�na�Q7៥H�'�_Zhm�Fr�k2�&�h�4 ݐF{R��CN�F:k|�E H��h�|����;�ӧ����G@ �����e��k���b�'󤀷�BY��� ����b��iɎ�O�5B"�v���EV�MU���n�d�o����oΒ鰡�v�q�5B*+6��=�ʹ�� |�����CĈM���G��x���0.���q����������]����x8�k�_��O꿩�����?b��#G|��\73��9����<b�,S�v���'�k�>(x i�C��Po�k�%�6� .����~���|s[��=�.J�%G��+�Mb�xn��
g����k��
�� 	5�)����������ݛ�=�?�{����-�~�1�Y��3���a���!�\ ���f���W�����z��+��~cֶ[��4��6i�zc֗֨V8����M�yU���N���4N�t�I���'���ط
��G�W4�q��F���6�ҮIbE���6�kh��9�/Q�E2��FV[%�ן֯����}���\��*����:VX㑘����<].�|I�U<��~&���)�}k�]��Gd��o�{S.+�WMеo�:�iK$I
������¡��ܙ�cq�}K��pi�:N襂���|h�N��$�s���`��Ϟ>�2:ռN�ᛅ�9>��j���{��S�����t6�Vt���v�w<'��M" #���Ɓs>#��[���l�u<�zW�G��V@s�f�A��Ԟ�s�8VpG������<3xo4�bN�Nj�
j�CP7n� L�W���j�H u��en���dx�C@K����Q�EI��z�\jMo9���^��u���S��1�pw+���YWpUb�]?��T3D��<SEy�}!��pq�ָ�[\k{7@;p=��}�F.lzט��7ڶ��Kd`��JV��K�ٙF:u���9[�C܃�,�%�bԬU%Q���m�0��"@09�t�tr}��>�˫U��1�?Z���ɪZ���l�X:�D�=t�%�F*�^g�*��T�X�i�+����tw� �t��`�_:x����n���$D�]lk7����M�^1 ��c���:��n�6��1_�k⏉��fm�"s�_E|#��ڬ��1'`O5k����B�b;UnRi�ɪY���\mcRdM��+��2��=�:�?ʽN�^_��nO�8�jl8�~j�H�[T�-�1�^s�X�B��$6q����� ���Wq⼮��KSz l�qؾ��u���a�,
�� �2���n���=+�5=݂�8!z��k��L�H2r{~�be�1A~q�����M�#�5�Zl��1�ֽW���ؑ@m���S=P��>���&��y�E1�U'�M��H�cx&����:��Ʀ�E|w�O��+� w�z�t�ҥ�}C�/�x�G[B��eQ���Ֆ]b�� �c�Φ�H��.�Xd���[�g���Rܻܛ�6kat��ʞ?*��M��4��v��1��|��e#�W�� �\?��V�	V, �1��96W*�1�#��f3��V�~^Ǳ���%��{HֿU~*�O�v����S![h ~��7�sC}?��Q!"!T���}�ғn�V�y�>����i���oˎ���^c�xK\)v:�W���@Q���#JͶ�w\U����ɪ���^��mWi9�fQ:(,x����K��=A�i�����ix�ǥ&ѱ��Rr�� J���c��G&��H��	���6�EC3u�֫���=�4�����{�֕���n\+�ݴ��gM�r�8��M���qҩ^m+���:�HA��OZ��!	&8�ւO�./R�68z�����$�i�o���0�H�q7&h]gp85�ڗ�}r�7�H�hy`»��#��%��|4�E��ݰc�?ҵ�0E���������z��?Z��K�u�J�V�y�H9�;�{��{�^�-Ơ���{��)E��J(��������u���������uoï�^w���B�>1x��D*�g�"�H�Y�I'���y��|Q{gu=��43\F�;���j/�����&I��K��egdݰ7C��>ݶ2��z��}�_q�{d~5��̃vtǥmfA�z���	��Mg������}�Cp�2c�=O� Z�t��6�C�|�zR�k��]]Wo�A�zε�d�fbw�ץu��+��TF�N�1#�)\gU�}*;�=�����gK����ε*��(�l8�����I�_<C�W�لN@����^6�/#��A�m���d�۹�g��xw��\ՄSK̒ 1�N}}k�_~�^���i�Ld�x�� ��zn9�+��œ��� �S�x�º��^���a36��<�J���<�nz?�/��f��j��q*�ɰ�����R\I�Lč�d��c����c�U�����Ն.n1�V��$
1޼�i6�����*�3�9��]xz����S�+#Ϯ,̛F@b{�sW���³<m��a�w�զEٵ#=�j4��N#*�|��q�]�V�����1u�H�"(�������@����(U���W�^i6MU��Ư����hТ�� ��>�/.�Y�O�m�!��v�`���l͂`b�z��x'��vSi�)~�G�Ĝc� �V�[A���n��t>�F��P8�GNvmC]n�����B�}lǪX7��0Hp+����쪲����~����?�`eh� mn�y6�uٌ^���|7ӯ$��C�;H��E^�<K�������^��"���l��#�d�X�����n�e�|��e&/3��d���5�蟲n��Gwّ��<�r`�\��� K�kV�{6|�� ��5�z����Vѕ��K�w�.y�h��ן6�+�9*��G�ߴ���u�f�;��ƕw9�.�v6	�p*��k��-oI��\8e�|aA�?�Wٿ���l<}��&7�m�\��#�[v� ι�/��\Y��Z���3�־Ѩ\���c��k�-k;�+1W8ێO�X.�$1�`����=����O��--��TE��@S��O_lׄ뭢M�}���#�� z�ӭ8˙\���>���i�m�l����`�3Rj�>���å�y)��q
�#�LW�o�� C��63�{�Hx����_8x���C�����@
O?OjkGaX��Oh`<� �q�?+6H�3���ںi��y�|�����Vd��}� OL���fb��UFy����A_|���SH�v4�p�(R9��$����#�"��ӯZ�3�d�����hgq��jn�<S�PX`��S��A�3�(��4�w �u╮�㜎}j�2?
 ��郷ڎZ�\L$�GLu���B��4 ��pNMN8����ҳ��ח��=1@��l[�9�oQ�R�����zg�w	���N�{
s9�f�$���})��}�HTmr(36H�מ�(��<��۵�A�Q��q�s�O�p{���� F8>�͛��jV��x�ޕ�5�wc�Zd����Wb��( 
���&|�xP:,!�g����^,���cw�TD�{�k������W��a�+��u>��E;���x<�M*�O�M����O`w0�=*D3q� ~��[ӜR2�)y�:�P�F�7g��NqMl�8�'��t��U�ۃH�6y&��󎇽/���$�(;��~� �J� ��R�-G ����� dc�
��h�8��K�q���Sw�q�ҝ�w�t��0K����9�)Gr:���`����N�;�8�=��4=B��4�Q���ݘ�#��=��Ab�ʨ��Jɵ�v���o��<:���F>��;�v�A�+�k��W;����3����G�Ӧx��9q��rIQ����Sќ��=)͕�y�I�0��~�'� *@5�����ˑ�Ɯps�E,q���m��q@hN�T�ퟥC����R��ÿ�]H�[��w��֣X�b2v�8�*�������}�_/l�Ι/\) ^3�?zQ��ړ��1�))v��J=h)y���h����3d��:�n�����A�l��TR/�	9���݌�<��� �͐	�sH�� O�ڛ�p��=�e��4�;qԓސ�sϽ7���qJ[^==1M� �>Ԁ= ?SI���U}��Vn�$���{¤��Qq�2<�8�}��"���{��[9���X^�A����T�a�f�5^��0Oo��f����o!���b!�L�H ��N�b��*O-���7J��$8F'>����~�,̬��x�09����L�&�����V ��^`�9�k7�u!���uc
9s#����w�'�J���?�a��*�_%ˡ�,�++点�b�a6���Q��b�<jD��W����ۈ��~��+����[[�%�-^�B8�������%���B7��=s^�-%Z�+!���Ը�Zf.�l���郊�/��P� ?�W�E��ʞ+��
/�T�r����N�z�T���l�{���λ������	=� _��y���Ukc������f#�)~�p9贇�}:S��׮j�ժ�)\�=0:��cn�/���o*[���c��S��f2�';�:����vs�o�j��m�)?Zz��2�-@�E����L� +��5mq��=�P�
.Ԝn��*�{�U�[M�~�x���y!�����VD���������6�s�@+��C�68��;~��xr=[�pG9���o�~��#<z�-���0i1����֮둋�>T�Kt*����2qK�6A�	�x���&[��`r>��~�{]4#d �V��m���«v�*duU؟wڂ���EP֊��#���V�ҽx��b4}8��2O ���]Jkp�sɮ�A[hɅ����mj4�t�Q�.N@�~�IL�#�clf�S=:��í�;	%O98���-ג[y��N�ҽN;��h��9�yֹumim%��b��?Z�.5 aH�p��= ��I8��;���D�`���8�z���c�0yu���tj���y7Ə*�`�ch9�X�3'�������l��H'�ԽE�ǐ���x�Y���>i���;T� ��h�l�H�^�� 
����e�,O��UO�K䵹�2;~��6W+�^Ӕ��w���\�ݬ���ǚ�c�������شQ���d��E{�=Z�<��<�����y��T�#��n�~=z�M�~ѣ���V�bp���wr|��y�����00?��O����a�ڼ���� Ħ�1��y�N��^]��n�=�cS`���'İ�����~\W�h�R��� �c>���j�X�G�y�d���lmOz�������m�Sh��W�jZ:�t�	���SU�m>0����y/�!�)��2i�����
�޺���XVk��� ����0�j�6��jo�Ⱥ�d���?���	�����:�����(��8��кǝf?�`�kz�;y5��E�f�9����09��=��u�eX��6:ׯ|��>_I�	�'�=J�/G![� �R�ᑸ�a�9��i�c�_������o!��5�²� ��~s�JQ�k,���?w��I�Ԥ�V�:�������+��a����Q򻋥���O��\`�{�����@�{��<u�E�"ݓ#���V�v���ƮR�$�݊w��\uj� ��h�2�{H�֐�7���_��~4�ۀ)��g�L	�{��΅;W&�9�8 g� �R2e��p9�l��5-����ޫ+t����f�~��ǅ@;�ֳ��`�K�OBO��H���N2���w�Y� nnB��=i��C�U��xP��.$��8���|�y��J�� Z�߄�M��[�Z��۷scW��H#�l�q[�O�=BM/�v�V�C�������z�8��8~�oÍ%�P������5�����爥��٬�!���ry�O~z��� �7�e���\��1V�1�S϶k��+|J��ڭ�����X��=�Z�[�(�<'��L�ֶ���u�<����U�ߊ�Դ9"�*��=*ni���Ha�8f17���g+6��<c��t~$���L�zu�W�.$���j֤7^;t�55��,��
���4ڨ[���+ G� A�)�����8�*�j�9*�=N�����w~��+^qJ��D�g �� ��y?u��g�}�,�p�;r0=��ŵ�1�0*��/�y��ո��0;d8ni̫�t���Q�u�09�_ƩnL�g�i|�xy�8����+u�İm�գ��~�6̏0 '�R?��
���q�x�^�?��� �VI63����-���<����_j6l�xU1ڬ�"�͐NҭXHU���-2��z�k�	n?��⤲Cn\{��GZ�(2QQH�`!x=�S���lm�}��}���dC
��n�z{WI$acQهҰ��V�Yq�z�[�z4��G<��F�V?�pB�܌�6�Z�;�0Z~���jk�C�v�{�=�e��P�枓��&Cw��U�'��;=B�B���Ic�`6�r� �Ǹ���h+����7�A�!�I=� 
���#�å��� 9���s�k�4� y�}�
��|e��K�����0!����Rk��C�k�i_&� ׌q^��]������<�\�E�����ך|?�	��ݳ���� ���Ӌ�N���<�↥ypҴ���X����(�L>$A3ac�8� tu�� �n�,n���+G�	�q'?���K�f�#�c�ԝ���*�NW�Q�3>�������1e۔���� ��1����2�@,~Ps�x�+�-^�/�[	� `	���g�W8��J��� "�]ޣ�
[��q�����������U�ػdcӎMV��F1[�̂e$n<��b���8�R�B#�֣U*����ך@L[�~`x��-ǐ�(�'�Ȩ��A?ҍ@�wn�s�z�;g4��+c�=�r'P2ǳ���DLW�A�8���7LՈW����c&r ǭ1��/JU�\�)�$=�U��dNMOp�T��CPd/`	�b&�|k���F��x���N�s�Ȧ��i��8��ʟ� ^)_����Nь��v��}��	�8)�����i# ������7Z�������A<��Mc�t�Hccc�$z�)$ d��X[}�N?Z�6C����@|݉�{S���p�j&bݲ3�M_����)շ�.g8�k�w�Rhr�3o�y
z��+�*�8����ּ�+uepSJ���*��!__ץ,�� 9=3V��x�W��T(��5���B���x�җ�NҀ��=��U���2�� ?6�>�r0�Hp[h��?g˒{t�֣\3����� *㑜�N�3I����"����:PP��>�J�#�s.ޔ�3�� E@��q����Q�Ҙ���K�O�KMbpG~�V�9t�EH��NMq�d�i ��~���5�Ҝ9��
W$��<�z}((���{9���S7��6�{�]�U��}�\��1��@�.#l�L�w�1�穧�rW��u����~��f?�������jF�)�Dq��LX{�õ �pr;g�ee���\q����lq�����s��}��n��Aڠ�^Iʷ��I��I/�'�*3�s����P^S#��>��s�J��{�P��0��bn'����8�jm
1F3N>� ΟJZV;�sM��n89�JG���0!*J��G�Ǔ�8��H�I��Nt��J�F��=�I�O�z��szT�� ��zi$�:PL~��Fx�q�y<���>���m���;@8�=)���S�F����-��Pá�8�ٕA#�.*1Ӷ)���z��N�\V@���[Z:.FA��ր;o
ڭƨ�q�=ORk�u��4����,zWΫ�M��1��0n*�2ե�F�4��i�M�=O�:���݌xJ�m[G���t�Ooƾd��M�2,�#!�?ά�x�V�b^���[�*�%��s�b�lf�%a��!�zDv�Dz��>^��������J�0>�� �T��=Jl+�ν0i\\�g��>Mc�yۑ�k�4��c�A.�qӞ|�%��w�3����� ����m�F�2����� ^��k�,��۹�s�����Bdc����[R>\y����Ӷňv��SѺװ�|���!��J�=%^f#p���^��N$�Pܞ� 簬���L�&�>��$��� ��� J�2Y����1��7`��Ws���$�5��˸�탏җp�ɤݻv=8�)��z�j�&8>���뫤��ʹ*�ߕv������2a��G�c��sǬ�=%ǈ����)E\�\W�xO��_b��e�H�q_���ʿ/�A� Ѝ}���;�61����ؠҥ�����i�b�Q]<��`��r:��%�Ď�I���@7�w�2}ι�o��麡���� ����qRۆ�h�w'�������c}����Z��84ci���Mp��wb�]x���"G8�����R#�� �&�%s���ZI��٫�MѸb1�{�r��x�{n�+�w��x�c+ `�� �wc#�R��#�7;�*�m�5�x�sk"8��1�&���DEV��k;ñ�h�B�N�����*��������X`{d��5c¶󙯤��y1��zPV���G�E u)���i�u��������z������+�����x ��X��S!np�z-���Z�a�*8�ڽ{A�h���*(^=+ϼ5�Ρ9�mu9n��^��H<��E46]C�'���85I6��"�x�Z���MW�,T�1���R+٦|��gB��n.!r��]Xp=zV_�&}�X���|�A���2eU��ה|Z��R�H�k�Q%���;�5x�.�k
�&�卸Ǡ�����b��F1��S��ݝ��m��<�
�o�>�����Wwҙr�{�%���� ٴ���cެ\a QӵU-�R3 ��(����w}��W�����p1ׯ�Y�*;���5�}�� g'��Ym�1q�{ύ-@�� rk�t�5.u���F�t�y�V���
�Z�6 ȯ�q�\���q5�F3_Ej��m.-���?Z�i�� D�A�֝�jg�WF97 �ɭ�9^o�W?Jʱ����"��}�����o(�}EC����F�}�\,~Km��w>�$����1���O���|��*���m5�qīǥa)9�D�&���P�W�f�qt�zWg�xe�dH�ްd�Ĩ��Ֆ��`��푸'��� J�Y�dg����	<q�DU�R��ɡ�UoM�߷Ҁ0�Pd�p@�|�N)ag��-���G�W����Y�¯n弼zP#��yf���of^���a�d��,d��[_	H�	a��)��Ij3���� ��Þ���A�9�ݫvO�
�P۔��s�jh�P��H�+�
`s�N��M9����z�F�����Ln.:xfT���'�;��� �>9N���=�e�5%��d~�zV�>&<�1#���+��L�Fc�L�6�y]��I�r��� *w� �ʹ��d`❐\�#m��"���m���
oO��5�܌���j����D%��Ehq�F_�q��kn$�{���<9-�co�Y�],�\j�� �(�'�:�;X�� }j��/�:o�#լ��.)w����	�ֺ��o/���0_ֽ�����]E���[���T'8Q�'��V?	��G��џ5�w�pi7Zg�|⡤ ��������瘔)$���O��W�7���4�ͼW�8�5a��J�c�_
�E�]ǀ�Yw�J�cW�/�r���N���>���WuN��>���Om�(u�zz�ϻv���j�x��¤��}sY���3�=WP���+�0�:����C��~'��p$�BEkZ\��288�;b�FĶsJ��7� �>���B�[�#j�:u�Dܫ�3���TH��1�� s۞?����$uZʿL�ޔ�,J�m�i�<25���'=�Z+��<���:�+	I1�q�Wm/~ʿ2�ڀ5㷒F���M��>bH7��T��̎~g)��
}G֘5��@wu=�S[�/���a �HII�{���sY+!��drpz�+Gìן���/�;z~u��W$���)|(�,b����N��
>b;~��-�F���ԑ�l]�X�zv�ċ��<���ڤ���q��5<�#n�V*���Y�I�2�FO|{U�&_��J�X���M�Á��4���N�'o^� �D�7�b��a,*
m�ˬ�����t9�:����!]����|�l�J�ݷ0�v�8�֧���`�=z�m1:� ��� �_�,�u�y��s�?�_y���M�M�H�9,��Z��������O庶F��Z|Sյ8�R��p6���+��RR��8	�MOP��>%/��:M��u�3{a�?2+����mlLS+�oS�� W��I�M��d�O$�k����z��Ԙ[��S{��ӧ�� Z��P���{�x�5�+��+*���8��� Z��{�n5�{p�7` <q�� �W����D�Ｆ���rb^8�~=k�n��W� Fb�F{��>������Z�q��`ف��� ��7hSP���Q#��}+뙯��	� ��6r{�y� ǿJ�CT��'8����7f��eV��x���������b[
1V�m�F�I� ���呲����C#�5*
����zg��R�{�Q.w�< �s��{�P̽p=���-��<�3)V����ށ��s��Tl�*b��9� �Ԓr�g��h�ϛ ��R�1�����ҟ���9� ����2�F?�=$+���r1�P{���Q�}��L	�Z��~U ���VX��TM\��Ɠ��H�ϡ��.J����0��E���p���ˀ��N����1F	=�aޘ�����5�ʞ#;y��jD�[��;Z@K��������w�ң��E1��&�����8隂_R���J�≣c��C��3�����o�iq�d�4��9{�*D ��Z�|~m��y�v��qT-|�
׆1rl=A#��V3�I�Wi���=��,��#��
�R2T��u�J��)n�@�n���c��@|6''���8>�^=����'�"����	6�ÜR� �c�A�i;����i��;
@*�ý9G8=;R���S۵2���E��nh���i �\9�G��@'$zR��4��h�������If�0�Z~��G-A~�v��;�'��Ry<�#��k�HA�Ǿi�#�׿�(�Ӯ:�n�'$d���֜�t����#�\rp~Q���O_�=�
B�={�@ch.�+ڕ�Ȝdq�NM6L0�ʊO,���@��2)�F+�9�ʓo���*�q�OjWY����B睹'�����lݞ�֍� ��4����q��V3�\z���"���r)yo�g��h2���"��:z��S�^�P l�!Yڥ~oЁA��R�j�,>��z�&��ҙez�j����)J����1��HGh&���'�f�����ٰ��g�=r�s��6X�>n��v�P�o_��5a�'�� ���� #/�;�Jg��~��^���j1�� ;���?�#}�q�zq�z��l�	����a)�߅@���{�T�(0nq��Z`U�Ӝ�j��ت���Z�F
����OK���J�i�,�0+���e��{Qt������JaFh�UUϧzѷ�V�^9�}�6?�`:��jû���:�������ƻ��sK6�^G<�� Zm�q�LE�UZ�f�w�KH�AL��������О��:T:����Rې�H��*=@	,�b���~���?�{�xB����Ln~1�t���j�6��^��]̞$�9Rn1XKs����?�T?٠2�]�,k��I������z���B��b�i>�Ҏ;{PV���2�{ו�h����<m8=;W��Nk�>2�7 �B�`�$|���C�0���bI�~��b,W����+��C��ęz��b3�&�@~�:i9��#J�c�mY-�`���W��^�����nq]/�b�8sg,q����L��#^1n�M3%������b�kwM�Ԕ��H�|A�HRM�.�������r}߭ ����7;U�޳5mZKXFHEo˯Xm1F���5���1ǐ�ܞ1�jWW�2mbǵy���a�k�>HA�u ���<'�Cu��P��PGz�:|Wח? �P1��b�EFE��.2A�6 ��=+��ۑyf���|��G��]���n� ����4d�'8�z�l�����r�4���9;rk��͜u�g��,���e#4���:��Wv���s� ֭�k��9�Do!��䢹m6���`�z�� _ҵ|9t�W=���JC�='N��%�؅+�~ ?�~���	��z�� �����<ז7�M��vi�J���m���DRpy?�z���HԮxs\Tt�x
ǁ3r1��?�u-���� 1�(���I>���i4{W,�p3Z�W'�ּ[�w��7�6Ս�l��!Z��>$�q�ϸ�g/+k˯<E�o)�`�c'��j/�~ok�jDȦf���}u��֑��"\�|�愍%%OC�7ǚ�������rx����]�Đ"4���<ԟ��eI*§�N����;y'��#[Y����1��' ~t��j����r-�a��e��cxP���щ��+u��i��HGϊ򿌊~�p:�W�C�W�|c]���q�Vύ<U��-ӕ��^!�k�''�$������U�+�+��+�ψ���/�$US�';z{R��By��{F��f��U*>\�r{�p25�\x��4UH*��*����)�1�i������;�yU�U?Z������ �_�+��uEw<���'��������y���fOX��%׏Z�_x�o//��+��Y*��7��x� �z�|���[|�� ��CM�md����C�u'�pC�c�S���ɘ�$8��;�WH�]#�x������� Ƿ���"�f_x��F��,��#�Ck�XJ���Rq���QqY�1���n�?�����0�Z�<o�݌{���W^476��
EY�D�����=*��0��rv���XW<���G�9;�{`�)��v��.v0�B)�X۴S�P��?ϥyl~2�o~jG���6���ǩj�oL �I�$�}x�Efy��"ƻ~��w����x�vV�j���%Yb�>p(�`��ઝ��A��i��V��!#Q�s�	��)�<P��-ܑY��0���/��J���0�m3/���m p:WC�<o(�$p���B�O���Ɠ�Eڣ��#?�HRG��!�Di�-��8�]^��;;{T+$��H��x���W���ˉ<��gdQ�B����I�W*wp�B�S�M�|��̿J��mm��\��z���m�S漼���=�O]��>;ǂ[j��������z6���Z�m6��i-��9��%��)�����W��kt� _;fO@H�^�nr˗��:�����+9b������;�lɮW���Ν�-[N:{��Ee�[ �N�^\�3�m���,Nzխ/A��5(������=*�}L��'���S|�`�]u��TK`���j���!6�v#a�2��T&��i����� �[}���xl5Rk_/�L��c�E8Q֝��y��AM�u��S/��v�Q�ɐSY$������� Q���� 'U��=)���ڤI��K�M�>^��W�)-�g�00��<)�9�H�웇9��4�.�S���5�����Ů<�UU$���KF/3��� �ҝ�,�`v���w���DlA��Ю��#-���ڈ�D��{�dk��wh Sʹ\r �}��5����>��3[�m��/S�U8u�2q��k9�����r	�b���|m���%��5���8�j���1� �lT�O���R�֪�����u���ٗ�~��U��;��z�FÑҡ���ܚ��̿�8!��%��������#9���A� u�}i�X��^>]ߕt�O�j�R�bq��wnz
���q��0��>�㱧a��Lʽ��ڵq� d�ӌzUk{�&l��v��6�ԯ'ҳl�9mR�7 |�?�z�t��>��I�]f�#F���/o-s:mȞs�O@��z�y�w>�&�`�[�f�&�����?t��A�r"��\�z�޼5�E��7Ÿd���/�᳼�;���b����B:�5�9r��b�<G㇁�m��{��F�6��GS^9s�����w$����#���]?�{}u|A-���Ф�G���G��\�1]j���y�0��sO�k�>������Q F�w6�>�q�W�Q��Բ0�?t�S_E��o�X���M�F@,�?1�ׁ��MN�q���o'�����T�sS'PF�Y �2+�W�f|���]��' c=뀌��HF:��*�e�VU�G���¤��s֙�F?�1�{�q�N�,��3� ⚤���zq�>�y㿵 3 ��ԋ�_J�7���1�*v���(���#��-�a�p>���7a-��;
�Yw1��� �HC$'�z�H�U�'p�$ ��TJCv�d�6EC��{T�����c p}��D��1��{Ч�)�>^��2� ���2=�z�>o��ڞ��9�ޣ��c�w�3A#�3Q������Rl�����*S#��#��Ioz� )���>4ڞ���g��P2=�d�1�N���q�S㏦yL�T�c���l�ny��H�+c�=m'�1Jz��*D$,W����+�s��)~U]m�G�=�Vl!����lz�V3&O���bO>�6�'8"��&'��4��㞽*D��������4��1�#'���v���?J@@G�Ꭴ�b��d<�!x�*2�X�0l�Ѱ`:��:P������ۻ�����Ȥ`z�z`>I7H�7 ��B���1#$��0��q@����ۜ�6�PsG4n��uiy��z�~��� �A ��w�n��4���}i�����A�zeĞe���1��L{�'��y�d8�p�^*?,�� ~9�1U�N��E�<�C�q���o͞�ݨ��#�4�m�S��� <��(9�H���9QN^=�qO�������FGZ��ޝ�3��(0ͷ�Jvz��he�0r���Q1���dv�		;I gڙ�+��9'��~�w��pU��9���v��s�8�֓w�z����Gb5�S!�z�� g�0[=i��y�۞)w� }zS������S��S��F{u���u���Ҍ��L��N9�FV�'�� �=X2�q�z�(^��� �K$$�9��9�~\g�b�������3P�ܾ��� ���e��)�FK�\S�
��w���	�{�����G��� �(Ns�ZT_�q� L�Y��?ҥ��[�Lw�����=�S:' �w4Ip�Z:I�0ǿJ��+�y�W���$6��@��w!�'��*�W��=��*�6� ��T|=s��b��$ͳ(U'�X�������zVż�4C��҂Xˆ���ڢ�^rx�����x�6����H���]|�9�� ,��c#5o����9�T��sAC��a�8�O�&��b8�� *}�^c1=	��� :/�;7g�8� ���!]��C���o���Mk��<��ּ+Mc��Z�_��� �QfNެ�>�L�2�꧳?K>��I��1��v�<�Ǟy�|$��� �@s�����٭�z�{u����?��9�Ґ�O��򏌋�Y��S�W��Z�M��c�p�R�#��2����C��ƾ��/��P;)��b���j�.�"�>3ׯ ~���+k����)�J�_�)���&O�\���W\��0;��8�����٬nݜ�,y���+ʼ��TϘ��M�ދ�F|�Q�.#�H��9�#�q�����}�:��S�@����)���Z���Ydn���BMƣq��Ǹ�G"���M.��_6X��
��60Dӕ��$d��^o�B�6��[g�z�^��5-b�ocY�:�������1��Y�fS�O��t�9��K�v�?��~joz��;y2��ȹ%��O��{��K=�烷%}+����}g�:�(ϯ'�+�|g�[ ���q��(��~��Z��`�̋�S����q=+?Z�[�)	�*��4#���O^�3��e%U�~b�O�� k_�����HCY����I�pS�o\�|#��vЇ�;��� �iއcj�}?k}��?0+��4v�@��Pz�x�"�)�[�pr�<*����������J1��ZЏM�0��ث+���� �a�;��ߏz i@��|�[���8a��w����Ď}s^3���O����׊�G���z�Zo�-�#�I�U<zW�V�Ŝ-��c�j�ұ���&�"�0�8�׿xo���[5W���5I�]JnN��^<�-�ѧ�YK7\�����E��m5"P~�"�����>�j�G��!��Hmd�����1�k�Do=���rT���ǔ��u�-s�P?�u����|�J���gR��5�:^���l��=H�R�k���/�i��Nk�s��o��y��9��V56��ڍ�hn29��U�Ƌ/�NG]��k�}H�pϸ��G����7��N#<q��|N�������Muo�V�Z.g�l|�a��i���zO�t!���Ŀ7N�����F�\ұ��7�D��m������ZM%>6��ھu�ik%��$`Jt#��kA׭��7Gbp�W;cTf\xvg�ny�*�a�tbw��~�\�i��qU�/���|���œ@N;㟥R�A�u`�J�o�� 1)�)�}k6O�p�L#�3 �8�k��R:�4�@*	�����cnH��H�H���\�m�GP�O�]���$�{6/h����pʟ�N>���5f ���b��x���#�8�T�/�^�2Ӄ���ǵ�C�]Σ�&nT�N0})[��Tlw�F\U(�`UwnQҦ��j�AA�����ټ:��e?�V_'���W9�x���[$���ߋ�S�(,���9ѳ6��>��{
T�Q�Y��z�A�Y4[�H���3ޯ�_�Sx�WB�����ʦ̫���}B���D�e��23Z3_Ok��Jm���z�X7^=��Rd��qޅq\ч����o�Օ�,SaH���+����m,� Wv끒�Һ�	��=SW�� 4��(�I#�斨i�G�RX6��g�:O�e8�=+�?x.,Q���u�g���Q�z�����Wr��������[��ͼ���#�AL�����g�s#�Ů!hYe_��z��}�����h�\z��'�W�� hYu�k��	�[þ�a�/n�I\��#��{`��^��8%�����/���:�:u彬7��r{�	���&���ƋQ#�T(����������.��Amv!حt*���}s��K�[/��3�r�m",�v�+���jg��&�e4��� ;�:՟�V��,����ⷦ�O��E�Ոǽ;^�ι���_J�KS����$s/\=��/<��s^��Η��ԜsU/�6}1]7��$6_jo��z��� �4#��Oi*����?�+���Y$c8���6�5�� ��*hc���d
�f������T#�'ṃoNi�����l�ׯ��g��R%��eR���ߥyχo- Y���q�~��5��1^9���\�m��.NS3�w|eF���� &�n����L�x�}�#I�����('ڭ6��g���5�N�O�gc��a��ϒ�ZD����p���s����X����ɏҸC#}�������
�`�C��^��X*�~Ƴ�����>+Ap����ҩ\�fS��8 �*��$�zp1R���z���?����8�c95%!�j�H����d!�����{T�0nH�C;W��P"��.2p	��]&蓒Î�+p�v��ys�X���ǥQh}���-�ִd�l8�"��R�`}�֬K&�3��V2;)�C�KP�[�ld��� ���]٤ʸ��t'��τ� �<u��X���ޠݑ�������u�/��&���x�#�6ch�'$g��x8�B��������;>X��������,�.m�z�+�ϋ�4�39�^=�~��/�I�iZ��-F[`ei�=��;�g�_'�n�w�u�%8��t�(�KS�^�1~"x�ͻ2��/\�=��|?qs���v����X���R�<�ry�<������F��W��$g��Qq�S�=OE�����H���Q��|��e7Z�v\rq��澮���c<~�`evS����?�|��Ĳ�g����]��X�:��Ʉ6�A��?
�"_��H=�n�g��G�Bz���er�P����ld�`s��8��7`6Fj̃��xc�J���n�%��`;�J��� ���#-F}?�E4J��'�4�#a�����lȪ:UXv�un���;8^{�+�|�1���r��J#�+g��B�q8�hP<��H���!�1qQ��L�#֤���9�Ӛ�/��8�*�N��g��j�d=H�S�##��C��ߞi�<.���Q�i��rp=i��`$����1��s��.�NO|Ҳ^N�Ml�����s��@9����/J��x�n�����u�D�x0�\�t=*�%�a�c|�v������ xI�I�"8�����\��9��ڣf���6GϠ$��Ĥ��~���!�_�屎�
���3��3Nϖ�$������6��j��T��p>�����OP\��� �J�Z�K�#��^1ҍ�q��D����C�FD����� ٵz+����z
y����A89�~�i m�>��")^�
T�T�GqMo�h'Ҙp;r(���҅�G
}��@��~t�U\��S��/\R�-��G+��)�=�y�4��P11Ӛ6�"����n�GҐ.�:A�x砦�x�H�ȩ|���W����S�r�zs�sL�ӹ�8�ښ,��v��
����,�����)�89?ϊc"����	<����
;�`��8�C@ۊ\qM�㸧/+��� Ni6���KJH_z E�Wʐ���)�G8��e��Wr��������9����R��An8��k���ޕj�ɞEiWf�r�6;u� ��Zz֣E1mi̌���Jy�\0���(#h9���E5�T����؟����gfv�-׏�ޕ.%W+��l�v������9�����?W%Q�(����U�������3�R�/�M�J	8��I�($)� �T��^���0i�T��Nq�SO�1�9���+a��s��,�c9�NO>ؤ `O_�r8�b��r{�t���ߎj'm���T�ͻ����*��'��S�|��r�лzqL������F��ץ��&���p���J ��R�AR��o l���ڢ�09#5h��ep\����o�hiq��1�ިpz���j���\���������Y�����T<�o����4� ����Q��V�$tG�9�+^|���۵c����ִ-�8B�=��e�eX�#�E����t�e�rIa��S��U�wS�@t5��|?$z�f��aJ�9�jK��rŇ��U�y aH��ūy2Ng�����#�9��m�7g�jMIr�~�d:llf pH$b���j��OfAKp~�ּSE]�n�H�^��]�^*� �w�ֱ��U=��O���Aaz����{��6y>¸/�-�M�q���z�y�O�l�1���e[�!��3�:rh_�֐�?�k�~3,g+���N��J��Ey7�O������ߦ*��>����|D|d#ܹ�-���3�f���������$�W ]6�: x���ȶ�`yg@y�Ъ���<>�����I� 
��|-t/�(a�/�}W�	a��e!UڮI�L:��U3��4�R<����e�F��+��4?��q&6j��&�M�F���zW��Br����\����c���{��LzƟ)`U���z�iv̸�UY�k�v��$�s���엒xQ�2�
����o�㽌���ԟ�_Kx����{J����)�4���C` ��~�)+�t�}5"P���>����-�c�aPyí%�)�W*���:�.����˨��#=>�C^���`>U�׶+AT�5��������MBݮ/�	���k��'��0��E��rh�E��g�FϽu�5�[���~t��|���3N�Sm�4�8#"�c��������-z�U�& 8�ג|N𼺴Q���W�&N+��&�䐿!I��ϒ[���ݥ�q$�ED߳�7_J�a��5A!T~Q<E�����j����m�y	>��/��+����Ҿ��ִ�۱3�� �k8�2�T��u��Viᯄ��>��_b��Ҟ�{[eH��5�?1*��G��#����B溱��n��<��B�N����^�2s\?ĨD�3�2�cSa#�x�4뫵$��p��_,|F���H�2I#���⯄P�H�Y�O=+��}�\�69 ⢛�"�ٷ�^MV��D �_IAcm��d6���H�N��H~���2I�<Kp[
G$�J<���>����+D� f����7ʟ �ּ*�������˰�\c��J� �ś�Lxo�� �W�+��y��k�;(9l3SX^4���ػ�����]C�����,}+�׿iiuH|�ŇB3UL/x�m��v���k��nu�cY7�;�<g=��j�]�ˍfG�@��sVwSڦT0��:WTS��7�Ϩ���ib)�*���K{��P>��M��"�ZB��x6���db�Yrr}�uc	D�W���8���b���Q����y$V�yy�?� �w���9t;��L�\�	}+Y�Nn�EyP��2?y�zWW��b�aTyWך�d��I�o�l眊��?�k#�$Wj��ɮW���"�˜��_�|	���?j��L�v}�l�kmO�5��^ �R9/�Ev	��i6�n I'�� _��_���"	Nྵ���ޑ"Ʊ�$��tSE�{V���,!��n�z{W����v3Dʈ��Y��F�c�=��d2)?7Ҽ�_/�.[я��k��4�#+�����4���=1֙���m�M=K�� �v�+έ�(�j��΍�9�� 
���Z���B�eL�ێ����sE-O�_	[D�h�Fp ���6���G��豷-�y� ��G
�s�Y2:���%\�����3t�s2�^	�Vݣ]ǧ֋!Y�W�%��X���V���^ռa�����*���d'Q��j�t�m�Ӟ=��� �����{�0M4�(Xa}1��]�he'g��^��|�t{y�"�@S�cV� ��3|;��7�w�����e;N�s���}�?�<1y<��C[}��V,n<��z����𿉴�>�����k�>IS�rp?CDۺDž�;�ˋ��9b�q�u3x��M��*<V7ËV��a۸� We�x]������H�S��K�v��We��z{�<��j��I����7�M��wFK��j� �0�W�BM�mi��N�t�� �Hш����d�cڧ�g�0{��@�w�Ep %GcUH]��G´�G3��/RMk}#0F;�Xf�]L۰��u�v�q��u�m��ds�Z�u	Y	#�9��
b3� ���7�=3V�y�%"���;�A�TX���Ϧ3T��kS�~���-�N��h6U[�ÞC���g�����ۙ�?�Uo��Ĥ�	�j��S??�7�
��������,#<���~B0g<�s32��}zև(n�L��M-��a(�;Q�s���&VVR���zjw��UPT�w:�+n��Ǡ�ށ�mŉR�1]-��km�PG�X6�L������>Ι�(ǿ��KSX؍q��q�R6g�W��?A�����:��H英����������$n��q��|Yw�#���χH�%�9
��?�ھf�q�O�x��(we��<�q_�_� g�ׯ��c���M��g�_9���S�#�0e**'�?#�� �Bbl(Pѯ u'�5��9�~ �&e��NNq����?�[ö�i�[�J�v�%U�0p@��|����-��˻�V@Wkg���ץiB�5&�-�uMR����)�@خ�W���Oj<�݌3ۊ�?�7.��em${�I
�$��C^=�L��Ϋ��w<��n8��<3�+�K���YʛQW��^��_,��R{�Y����������~�}�/�;�9ʟ�z�(� 
��Ve�ԕ����=Ltf�����ӑ�ҳ�79�=���Ze�X���T%����?w� �[�*��F�I��F�o����\s� ?����Lld�{ԅ�t9������ �]��~x��Q��P��ޟ�HDl�I9�ވ$m�����>D�׷j5�8���@đñ=*5?1���RH�ؤ�6��Ͽ�@���9ʜ�xg��S�9���	���A�qӭ�|����PLy<�޹���+�s�SJ�|�}i���?�zE����E�q�Ts.�\q�� *@Jц\��MB����z��eʟ������\�FsH��O=)�0ǩ ��քʱ}� �T�N>��1@ʫ��7��qM_�����  E��	$�v�6��)c�7���SL�v�:Z@K�|����ս1�y�:�X��%���c��	��5H
3&f~s��֘��#����J�VwS�z��j6�pW��Rz7>��)��I�#����v�BOJ���Q�pA�4 �`�;;ҫ��7?«�QN�Ϙ0���( -�� ����R��s���;�R��Q��~�#\�q@x}�Lj�d�FGC����?Z�����'^{��C��}�֗�>� �4.��L�,޾����=�S�TҔ��C�0m�t�R��+��i���=)O8�j
Н��.�A��99�,��B��S��0�;����~�q��P���I�l,�&����{�sLl����� 9r��� w�*�q�R2���P3�b��qϽ#�� �B�^�#}�@�z�@���y�)F�@#�8�n9\��s�vI�8`� m-�84���dg��V�0���n���U��đ�N6��@	�k0���zR��'>�2��ʑ�� l��i�G'(+�z�4��F{R4gU�(
pqY��q����C��]�#\��>��fwN�=i̿xO�L��8��sL�g����Irq��}($���f^x�t:~��X�c�4ym�$�A�N9�MQ��keۑ֘WV&�FRH<���͑�;q[:���8=�V3}�t��Xپl�����'�H��)�����B7�s�Q��&�8݁�s�>�� ݼ9�iQ6�{f��p{�e�l��P�/M�qV��m�l�;v(���\��[wn ��Z���ڴ�3��>��8�ֵ�XVln� 65�_.6��?ƩD�L��ҭk2�����������;y-�#D�71�#���S��rj�K �c�Pmܤ�C���	4��Ԛr��(>���^���z0留oI�I-�cz属���|=m>�@�(\�9�k�{=:�C��7.�%���%�q�׎x�P���v��W�s�u�kš��)����Q<�լ.���<�ҌS�Һ�YĪFx#�\td�}����s�W<�Õ�Sh��I��
-U�����]|А95d<:�����װ�(e_Xdm�g��J�� /�� �5��� 	E��l{u�`�#���Y���i�ɏs^��;����� d� �z����5�,�3|�k�;�1��wlf�F4��ɠ�����W�#D}R� �����n�Ŋ](F����M�.�����nV��>�?:�'��,�a˳·�k�W��1��,<Յ�`EeU��:�J�39{>]b�� ~f��+��H�aCU�w4����HD
/{~t��%�'4�w�нzR�P��t�!V���zR`��@�h�?0��Wv0]BS��T��qғv�⁜�Ɠ�;�ؤ9��44,8�)!K�7�t6�q��sX�"���ʔ�Ė�����G�Z%̒����V�4� /zĿx�q��d�b��<
�����4 �!0ZƇoʠ
]��S�q���l� /(��4v��(�"��`kZY�f#��o���P�����z	<��®�m���ǳ�*�5K��x�e�m��i���9��8��H�|�N������=�D���'�P��� �P�Jѫ�W��������5�m`�����i6^[(�AZ����TG�u�*(\?�b~�;�3]�lCq\W�?����s��q��w⾺mg����G�_%���֦bH;�}c�kF2�O&����|cǪ�N\� �*)$��o�W�w:���tfN�5�x��/��t������ ��mS�v�:%0x�� ��4�4�B?.2�v8��ne^\���  O�Y���_�e���գ��3�8��~�f�P�wm)�4�`Kw�?ֹټ�^<�
��3U�%S[X��
�	���\L�7z��>,v��#�k�k�&BG�A�#��U�º�e�Q�g�gǲx6X�謶�n*G~���+�i$�d`pj���k��2���8���^��E���%jg��SQ*�z$yv�����aJ}kZ��UTaU{t�S�����K`��u�3�u�K�_j�܃��j�����l�U���Vh��6~^p+sN����X����sI� 	S�8?Z����#8����98��\b��'�.7�=G��E���*[�z��c�g
���� ר>ĒI�ֹ#U��٫cygw$��bc'w��g�?E�Q*����y��ň�W8Ew|%?�4ٙ�(�A�Z���}NZ�E���6���X��NH���ʯ�����x�8$(I 8�l~u�|4�&��=��Jİ<7NzՏ�?Mc�Vĸ(%���lsiq>2|R�K�d(�_����^c�� �����6��Q�� �O�ks���(���
��Xʿs�_@�(��h~�<���  y�=@떴�K���Z����~��D�<c$c�Ҽ��W7:��VW��p�������W�wPIF}?���o4�� �������	R8��Bk�ToC��u��M�S#K��B��RG��8�śz�)��#�n�rB��5�G�A<Ճz��<�C�i��c�0FU���8�zR$�<���l�W���<S�H��݅��-؅f��������l����(,�h������#�3�O�,n
�<���z	h��濍>x��ޟ�cz�F6�O�=G�Z���ZԾ!4kx�b������ ��s�[����"i��"����#���?:�o�4ռgks~��e��p*ԃ��Q�[�j`�ɯ���k����|���-u	mdF��]���\��f4��_��� *��Y�.��-R�E��.1�"�^���_�4��Z2s�ڴ���G��ˌ��g���K[�9n	�����E��9�Y\���۱�ZVmb��eV���bk�>[|+goV#��w��&9�|�QGY������<�.�sV-��w-��Vk��C!?�B�g�c�Uۃl����UkQ�zs@H���5F�"�����*췑@�`�G���hO-��'�|/�6��c��1��������v`�x�t?$A�y� ÐO�+l1�1�r��1��ed�W��B�2?:��5�Z���6v��s��)n��S�{v ����26ebO8�OZCD�!U�N�j&a!�pry��֤3.�G<sU����ɤZC�Խ�q������ī
�p{�+��!�U�+�:dc?ֻ9��Ɩx����9����&:�d�OJ�Hz���zTX%��a��§���ܜ��RѲgY�F�-'�p��~�_��+�����f�-�V�����g���]R�J�P�!�?CO�������%#�U'�1�ּ���ާ���%���#\x�I�k˗x́�g$t�9�W�.�����$}�}�ǒ�A��W��j�֚���YN?��ק|%�n�{��;G����	��F<�C����|^�Λ�k)<����2:���߽xϊ�tF�o�?���ϵ{W���A�>s��>��ך<�m���99%INy�$j�=w��y?O������������2��n������`������xm��/$b2I ���-͑�k�h��w˃t�Ҍ��w�7�v�x�v���8�����X���(U�#��k�L@J��z�?'�Ʀ�z�w�Q$�ずG�=�P[ʖO���#�TMG뎾��=�JHC$o-y�=���Q���)�(|����Ԇ�w�@��_�D�Us���f��
�<(�TP2WE#��������J�T�*�g�Cc����0%����w�{S� ��z"����g�Sf������T2dd��1O\c�G�H��J���"�eo�Q�����M�9�<�2L+cF>ԀU]��|�M�v�?ԉ��ޟ�G0!Nzs@�#��w���*�zn ׽��Ҁ�[�S�b6囡o݃���qNC��9�#�@d��?w?CW��^�#��=~�Q���q��_�Ȏ��A�=@��S�C��������LU�֥��^H�$���4����4��r[c�H�/'�4}��$�ғ���H�^�g�?�=[,pq�O��2�2qC��� �mv�u4�,+���]�>����ܧ�í0���pOQ�R�{S�8���F`�v�7R�$x����8H8��ϭ=
E-��Jw�J�f#�*6�� �=H��'�*�<@��A����r��s�7�v��	�|���Q� 1���I�OQN�\�$PY$�zm�py�j��=�I�[��w�\n$O�0#U!K�����B��;�}�þiʻ}=�� 1T������� p�9���u�j]�� �;�ڏ�N��9ϿjC��{� E�H2G��"��nO�F����F��sP�\I4xs�qQm��3ӵ5���ZV��q�@����qHX�8��^���@;r�4�.�����V�"P��y��v��F���'�j�x9�Ґh;�1�y��L��?�I��RN8zvZd1�B���$��O
�1i:�2��ƭ׵f��>�3L�=��� ��kZUƞ�[��O#�����bN�I��:�OY
��懨��U�u�=)�gV�}j7m͓�hy<�m�W#n���1�>��#3���H�H����&����)�B�$������Q���@~x�Ҏ;�t��y�#�>�4���9�	a����XdS�J��U[X���W�� �a��;�LFB����� ���8�&;2���[~'p��H�my��<rpj��� �w\�X�e¨��1����*�#9
v���z����b:��9� �k�~����o���Jѱ�?v����,tQ�$�ϲ����=.ԣ��޸���f���%;��8
:җN��� �RU�rC��k�?�Ey݈��p��O	D����Xb��<�N8�r6�<���=i��j�,���3���_��1�u�^�8�O2O�ܻn��RGu��
2q�j8[���bO�R\)�1��ҴFF߆��i�b�bzz���,�C	$^��*�~]Qm�&X� �.{�U�xc��D�1�����5��֦��>��?���``�p��^�3+ #�?*����H�!�`
�2k��'��V�ە�֔d}���w֛���ީ��	_�}���g�Z�E��p{����mb��\�\����@_ �sCd�� ���H ݍ�?������OƝ�w�d��n�Yq�ҝz۳/�EЍ0�����&��^�O����6�x���� �(�8�Z�� ��߮�K� 	 ��#ۥD�~����&:�j�� ��߻=�� �f8��IA��r�e����2���/�mۍ�.f�v��Mϧ?J�>%�8�?Z�pg���}(�3U��P2���"����4�I�ןq�.���fn(ݻ ��Y�V� ��s���(?���Afj�+���ך�� ���}q�� �I-�}���p�5�7lR�,����I����H|In�n�����ޅ%GJ�� ��ߡu�;�+r�8��Y���� 
RĞ+#�V���p��b����=?
�� 	��YO�M��6����?C�1>�k��#^$v7����/��EϮk��_�K�nD;��y��!��>~��s4�@�k�O��z_Mٯ��U��}GO�gR=��� ���A�yB���N���{L~���?��%��W��֑��ElN����w�ʺ(��������H�ik�)�����5ѱ�J�K�g��ᅱ*G-�>��כ�F�D�'�He_��z��W��K��O�Ť *F��������~ ��m��}�� �4�(�&Ϡ-|e��Ʋ� �Ң��:Ŝ�A���9�Y�W�c�ҡKw���ӊ��Y/�4WY�?i�2��-x�7?ť��]��_��}k��q�ͼA���g�\c�;�'�m-~)C'ʥgC�����W�g�M?M��޻y��sN1�sn�C�~�����mB8����� Z��_���]�c��� �]���5i��|�7Vf0�,����լ�!*���=��ur�*Ћ�e�|��� �S�$�n?Z��c�\����&�y\����_�m�k59�8�6��=
{�P��~|7�:I<�͎\���Um]�79��j�P��#dc�rr���r�0���2��V��״����
�- �Qǧ���&��/��m=>���컣�Y�;7��y�.~�3�lW�GDy����������I  H���W#�O���YE)bE�=0I�������W9}�܁�G?����t�l�<�9<tl���R��*1�����DjVV�5�D�v�[����}a�O�� ¶�����b�}���}�[{��b��}���׫�%�T>��y���n�y�+�]'x����>-7M�E� �ש�|%��/�.KI�E�_�ӝ������"֠�þ���̥"P@���+��8o���?1����WM�l������f�m�NU�H���]~��~5�� 
do�P��tW{�1'�V�1��Ԗ�S�v8���0�j�[��HG�T�����*3���c[͚e�n�;v��y���\������� *�V]*�GFۆ�Wm9_qN*�֞2�#m��A�hPG�p����pTJ���,c�<�#��L8�rG?ֹτ����ܑG�90���p+����3��R�����ؠ%��0	������2Qh��F�F�� ʒT�����i�J���Ԛ3�=k!���u
jb��G�VT����jd-�l������c�� ���3�Ğ�Փ'��'�ԬO�}@�+�c�����ry�6��cv���݂NӞy��2H�r�o�jB�$8��Գc���9��ch���TX��R���q�9����V p)�&����}h[�[C�7���o�)9Y��x��-d�\�Ğ�Տɷ���, ��!�?�E�\�'<c�{��~q���H�2#'=�7|�d�_z�p���5g(��ӥU�~v ���5>�?�ԗQ����"�M~\�'<��Hs����~b�0>���͜��U�b��R�vFO�zߺ�U#-�|V�9�s���.�=8�-�Kr�'t-8��x������(#�3~C�C�X��{I>��0܂߁���,��-������t�o�J��bq�$�]f���N@�=�r�l�_LR���z~U����L�N�J����x�༕�J�߇k�^[���.����;��\-�tPF����>��!��w�\�g�q޹�=t�1�AUv���~nrG�^.B���g�a�ۊ����^[�Wy��NNq�����V�t����I�Tu��c՛��|?��MN>�<�z���z׉����Ns��׷x"�Z�r�!բ ��^%�!]ZU,p�s��DV��uB��͌������L2��kB4V��8L���n���d �n�#� �Z܆3����� ���.}���Q��_���C��{ү���F��C1�])��/��u�O_�}q�4!������Ke�NM�vNq�#P�N~j`:O�P!��9�;Չ��E������jC-�<��`��a���T�'��J������0�F��f�L�A���4��<q@�@�2�?�5�f���O9\�׵5�z`�P��Tq�Me�;�2?RF�(���p:w�zLB���%�aޣ����	���������zJC!�Fr~���R�����.Ӎ��;H����G�,�,H#�*ͨı� �8�����1���:� ��̌�ۀ~����I�L��^��A����=?Z��m��/=jޒDW/���������|�?Ι� -B���bFs�����0����� W+�;zqO��\c��߱���3Rc�[!r3�=)F���ʠcsNV;�c�`��"��<jR����jg,����) �6����;��sv�A����n��8gh��1��l�rO$���y���<�Z��1Lc ��qB���x���.T��@�ϧ5"�$�cc!�K�Nx#�d� �2�p�<{�O����29
[�Rǅ<�����c�6�7��ښP���֕�n�� v�9��� ^��:7� ��F�2I>��������p'^��}����K�p|g �ր��\���>� w�;��6�q@��Q�C1$��� P�Sj���օ��t=(|�·�4�BXϾ?�4ܶz��#R�r@��ր��랆����qK�1�?{�4�� � �OzD�7�mh�I`40�:S��s� �l60q� �`U�
��F�1����?A�sA"?�1�c(�#���^�c��PYF�z��01=i������})�k?�M݌�۵+t�M᳁����.��5a����*M��G SJ��@8�l�~�����ϯJ�?@A���� 1��v��H>� Jw9���OzvӴsאq� ,w^®*���;I�栂-��^���xA�Zנ��b&�@�<�S��o$?�d"2�F���iGL�^���C��;c�Z�D�� 7r1�5�z�<FK~&�7GM���"�0}���4ۅ$l+�aI�u����Pɴ��n{z��� -SCI�Q����Z���c�浚;Џ¤���uʌ�S��]� �+4��
�5sᮓ�y刳W��M�\+e����}�c�r�*{t��u��� پzF�6�Q�g�\e��kK��u
7c������i��O�e�bq����щ���_NM�~����dg�SY�	4�f��Ё���G�Z��NO���9b�.ǧ5���/���Bw)�*x~�-�%�������5$t� ������T��O�Nk�~*h�w�IB�s���'�~��#uUT�^+���ƈn��U[r.P���D�^F?�u�m~�&�H� 3�A��A��y�۬a{s�|���[]�R�����]M� ���Pҩc��q�ݝ|ܧБ�|�W��}s��#��ӓ�r?�	�|��0&P9������-��BH�X`�ME��v=�����ɱ4�s�\UO�ild>�>$x�m�m�I3?Np�<��p�������楦Td������ُ�@>������J[�j�"�o]��C� 	&��eoΧR�����4��3(�S���f�q��+��H/wq+�� �2mj�N|��'���\�G��~Ұ1m��?QN����1��3��~��Z���]7���5��s\m�����Z�&.t}�'�˟���� �ҧ�	??39ϮM|ֺ�{X\�֡�Y]�<��@8����v>�� ���1&N{�<�r~�����H����C[�;��Fk�l�O�9���
k����u���pF}i��Ą#9��+�k_[�-0Ϧx�u'�&V�HY���V��g�<���O�����9��T���.f���W̚��`T!&���Z.�C�M���8��5?#��h+�n�ݾ�]����2 �ã(?ʾ^]r ��9�Mu�M�����*��G"�(������2^Y)�:�[/��YP�В���'���ڼs�4�� }7�D�Aڪ�My��[{[�w����t�w�Zg������`ߍC7�;�� ��ǡ��ƶiq��`j9<[l�q>�=�I�2>�����,�-/�T`��.gb�w~0k��{�QJ��s��F��"�C��rpkE՘�]�D\p|ϗ�5/�4l��Ĝ}zW���h������B�]�@H�ޭój�U� �J:�t��W��r1�~f�AMf93�2�SV���|��Ԩ���G���Ns�@Q� �E\]D�I��Q� ��H|c��G��[CG#+�yi�W����q:��Cf�����Hѥe$������ ��C�9B�y�^�a�Nc�[#4��e'�}��cN��e]��zgڿ;?i/C�j�I�<}k��G�6�j���^�=ZmPy�$��Mm�%���˯j	";�2:W��7�	m��<�wz�b��9㸪/�p@����~e����9����š�#,�x�'�mp_�o4uۜ��ԑ�oTԈ�m�aۊK��*<��\��v���}���|x�%�Er�8x�G�O��Kr���N|�c��1�fH���5,��<3��j�MKDf�ֶ6��]^kͨob��zb��.�}=�2�
����zٌ�$�J� �g +@Կq�%�4�_xzS�;F3�������]�L���9"�Nh��9k�~��[u���i�5�u܉&�8�k���n���;wa:���='d�RL`�`��K�.���G���9�s��=ÈW��(g��YN)������JmIn�����i�jG���}w�xzXT3ڒ�s��ױ���b�@��<����y����N�Q�lP2�z���F�u�!��ddoU�s��5�3kZlq��q�����ޗ�٭��JF�\b�cR��yGƿ�������2nڋ�oָ��%�l|Q��4l���ܜ���?¾�����j�fC$l�T��5�	�9�hv��[���w�[yH�!�q��+盻�w����ګ��CvZ����4���̬��6�m����V� �mjF��1'���kI�I"!��Z?x����f٥�q�μ�?�_���W�wMp�/]�z�6�m��$�Np:Vv��3X�%�[ȭ' ð�jAE\�RW�G�_-�z8q����=O^���5��C���� +��5�[�w��R��\6�?��{�����K�� :����(B?u�cc(���nE&�@G�s��{쵬�@�x��T۸;�յ69�h��d��8�a���&����d�i:�qҵ1����@"��H�0a��T�09*:�z �F��sO0?����+���
2?�v����Eg<g�J@iZ�^��D�А��8�5����3+뻱���Z��[���c�k��7��s<H�����>����-�e�/3�UU��9�'�j�-��T��b�{�]6V�֝�D�m`1��jmŔ��S��� girsۊ}��u�;F^29�N*�"���71�#��̳+:0��u���V�Cneװ�;V��<Ě�� mRG�qj��K��W��r
��u��Q+ap	�]�m���#�i2WӁ�������׹M�����}&3�c�gҥ^c���׊N8��.0�g�ZX�>���l�����,@��H��f� �.�EV�3׎:Ү2p0zS�3��T����Ք�8�*M���nŜ���kv�e��8�ci�ZLr;�h�G'��;V�
�ԋ��9$���D�����q��r1�j���'ٱ��c$�N�95%�sړ*T�N8������9�d�uH�Y
2��C\t0���8��z�*�}6_��C��ncI������n4{�@J�,1X�Fz����3^[,�(X�5���ue�߇�������5�v{��>K���+�OZ�y2������5m.�I� RZ0�����v,���jNcR#�zq��6���������V2ܤ����U�C��<.9S�G�5��ԫw�JS7�3��׺x�M�O���I�>�����j����f�<R��
��Q��ʻ_ނy� 9�TQ��q��ҳoH�<�8�&'^sQ�x�:���X�4r��(���w;M7>��<�z�@B�*A��z�ˎ��MT��'�K
�N0=�D��*s�%��]�gJ`8���j-�2����$ny;h��qHC�UW�ӎ��y[/j�TH�����$�ئ1��as������Zr���o���hE��g�<�e�c֘�G$�R��q���\󓚏q�N��
�1Lb`�� �s���Q��`�1韥<)�_Zkc���������!s�;�HT0�����i텐�9ґX� ����R8���O�������W�>�)�z���H�9��ի�}�$�RT�ڪ���#�\��+x�<Ƙ�����Z)#��W�v0j֬�V� ꣀMU�n������F76H;G�Ԋ�?t���� ��Ԁ�>��hEP�w�z�&ߗu�9�$q��X�9��@ǘq���Q�'��u�J�!GQ��o���`v`�>_zx^�}�����@;��=� ����I�?փ���ӎGQǽQC9���ӕ���zV�G��"���2Ǯlyc��U<�l��v����V!�?Ze��ѷ{qO��Q���=)ˍ��H�h㱦�/�:jM�ia@sN^�v�.��iKn�g`�d��>����L��:T�)*W ���?/jkH8l���b�x=�����v0q���?6�q���,q��X���4�W8?^)�n�VU�u���ǜ�@㜓��Jcc ����4m,݇�/�=A����i�� }})ۇq��n��ҁX6��O���+0N;Rn�9�-�s�	���C�?�j>�����㞙�A Ƿ���"���9ϭ��c��e}��.���4��I���;i���lj�T��Of��c�3�>�4�7nrT�)ʧ�H�?�M_��u���b~^�Z@9�\?kG��4���_�M��P�R��G^��>20?E���g�O� �� �b�p��[ZN��5�O$;X�0n%�@#�VU7��<��*�[Q|[�+��K6�(1��CKO3�����U��yjɐ[��֖���I�敆w���x��t����_Pj�1M/��M���3�rpq_6x5�Ė�!�@�a^��O��T?|�C���#��kT��������x�;�[SR�,[�9�:u�����9״im��w�8c�g�k�>���m.�1�C����	�R��R���C(d��lp��
7s��~��Nm���{��7����h��ھb�u�sI�So�&��P:�緵}���K��"H0
�遜���o��;\��i"B�C�Wk]O=K���ꗺňv�t r�ۊ�>"x�_7�/v�J��Z���=�GU�U	$��ş[x�^[;H���ܠ�������>U��5�ŷ��yu���t�����n(�;��}�������������cz+�}?�r�G��t�C����׶r*����$�,���I~�s_u/��;�bR'�*�|�H�������ޗ�'�2Z�W��Z7��ӌ֓kZ��1���q��> |/������s�'j�%$q��̫�UFW!�f���(�#m�ִ#�f�" ���c�`�1gs�Bg���*��I�7[�Z���nŕ�g����#{�]��{�A�o�2�;O��?WU�E.����t�èƭ�}�^Uzӎ��N/s��~�È�=��?�E� V���u����8�N�j���8ay �׊���D����c�φ�O�iYw���8�o��7.�s��
�����X�C.2xO��t[��4ؤ����Gc���s��?ƭ[�<*�[�aU�ˑ����*ݪ�'��\��X7W,���	=�i����h�d-�J�O���H��O8⽋�~y9dL �_j�R����g����@�!n�Wa7��skf.$,&u�"����=���E�;Oq�^�7�<��}��.qY)_V7�V>_����2��T�\�<�x]��E!���5���_h����!Ͻp���Y�yV��F�����֥Tkr���~^4�p�s&=�Z��xt�ׯJ�<[��|?�\��²1q�+����s���us9Ǖ�Қ�E^]�������I�<��(^��e�4�@�x��Q
�^e�0Ho�ZV~��l*I������G�-6�t?�{'�|;f� gޱ��<�E�;��)%=�4�_��g��8���^��)1�[�+�ԾX_i��N���5��)������}��,sn�>�k2�᱐p��^��W���iѬ��qmc�z��E�o�V��~���g$n�ZLe�\SdW? $� ZM�p銍n���>� ��U9##�MY���� ,}y��m��cE �n��ֻ��ul��".H�>٬܊H�|p��9~��n�!
�>k�4U�� ё�~b?�W��h�dV�U�F+)I��|7�x��H!Îi�o��HT�=��xoO��`��3�����7��o�����Q�p�<��b���޳.ː1V�o�߷? �M��E��/�l�33�,%W�Nz��� ��x��+��-	9
G��y���I|M�[;5Wn[���޿H��2�¾�3���׉�b5���Q��g)��
��mW�c `W�߇�sjFU3� y�^���Z�C�($
��\�Ͼ�����t���;�g�#n��+ɥ
�5l�RQG�zO쿧i��k�W�G������_,�m��M�����*O�����)i�ڃ�n�ce����?�+Ş��<W�4>d�q�r��סNN���/y�G�u��e�[�J���U�oa�x�p���%^����s��]*���ܞ����X��O������S֯ۼ�ad��ǡ�j�� ���=+��v��ǈ,-��'�[��	���t�g�����KV�����a�~������ap^��V�k�h�1�p��c �+A��}o#ȌJk����.�ѷ�	Ӿ���p�+�d�	�x�	e��a�>^I�1\e�ŭoTX-|͐��ـy��� �u[+��;^���A��5.O�:iG�s��g��YIs-��c�FI~ *���TԴ�A�'f! �x9�~�|w�ѿ����,�� **��9'ҿ~=�Ik����L���R�Q�̟���Z���"�=���n>�~c#�l��q��-��9�)ճ�We��:�ח�6�،��y����O�p�(�d�fl�����ܴm�F29���h\�/.��H���s�O�g�Һ�������Fb��Y��+��̛7s�H&�?����C�\��� *¯�tQ��կ��f�ö@���}�z�(V"������_��Ȥ��[��q^�#nr}Ms��_�6�2�4닂܁�im΢�h�� �iؓ��R��LW�)��zW�͕��=�ֽ�U�M�q���7���h=ǯ���7w�'�J�E�7��Z�V+�`��BH���ǭ;�F)�0(���<zz���*�pNzg��}p)_�a������6��³��Z�#�^�����𩙢"9	#�_Z����v�8S�<V�|V֖ŭ"��m�e�vV�����ڄ�Z�6��@��j���4���:W'�i&��2F�lrI�kB-aQ@f�����j�	� =��5��-o��IJ��r?:�X�+t�#>�}�9��J��c�&*;E@�����"������b}�@�v�
��#�ӵ�wZԞI����V�����_r9��ϯ��z� �a����X�F����z�� �֗���A��M�# ���J�T�FKk�S�<Ge&�y�Y�PZ�<*�{ ?ƹ����J����h:��p?yz���p~��F�6*ïC^�ISW?;Ƶ��ݡ� z�O'�b��sڤ���F�
��<�����9�c�Oʟ��d��8'\��f�s���1����M�9�@��ʑ�ڮ�h[s�n獹�\���r�v�{s�>SD��
�v����8�啍�g�w�p[�� p��x��E��� ���U�j~d6��J�pv`F�@�=�M${0H����Ս5Ws1��zf�R /v$�pMfٺ�����4�!"9H�+��+v�I#q������]H��j�bV���#����95�V��L�u�]Ԟe�����׻�cZ>[_�O3���ȇ�������Э�A�}5��ƫ���3�"У������)�PB��'��q�VG��S�O�D�4�<��U1�\W�G������)h���3�_Xx�N�Hq8X��
x9�'֯�A�x�U��^i2��/��͎�|$F�!�'�����׆�rYk�Г���$q�'�+����F����W-ǯ5�gĨE��f
pwrY��I?�?�%b����e��ӭd�c���A[r|�`c#�b�5&��G8�a�Vڃ���u✿���n:S9���AւG�ɥ��3L^�\S�ڰ�dc!-�8_�J� 5xe=�^je]��j ����)C8�(�x�S�PzSFm�P�7���I#0����{u�ZV��zB,��H�v�����RB6�O��$
["�G&� �q�N�G�B�8� �qI�+��t�?62),�\d�)���N��{�����G�&��s�jI0�
pG4��6?/~�HO�ہ�O���� �ӥ�j�O=�Ҁ!Y�q� {��<2�zR`��1H� ��i 1�pN���ӿ<f�Ĳ� �jXb��8�Lf�7�89��
6iCp������2�k��}��uI$�v�D���p3�5HO_P��)?Ω�Kn�z�ɫ:���w�<`�e�V^23�F*���0��S�9
8�1�UP��#�S��^)���!��$f�=;��<�C���2u9�ڝ��)�s� b1�g�t�.	1'�S���D{8��
���q���� �G׭�9$�Af���AB���5"�w`|�� ���ՋY����?QPmیә�	A��Lo�3��˷���Tʮ6��wL`��C�Eh����ջap�=���0zZ���� �0�e1�����J��Gzfe��Y�� :Ԍ�,7d/�~q���ѻn#>��c;�qF�U;�Tm�	ݏ�>�����$��x��J�I>��K�� ���ϭ����:�M��1ۧJkFW$��9�W��@�E��0>�ʦa�pO)a�9㷯֟4k�X��@�UIݒI�ޢ�h�=��W�)}@���P��X�Q��<w4�����$�h$c}�GzF.0N+�O�I�6O��"C�q��JE#v1��+ Ow���i�]����y�4�S�<��Sy�i2y�~M 3�^*M܎��&=�@�˜�V^q�Rs�Z{G��N����+]\6r:p�}(>N�v�?�b��C߽/n[֓g�;})�ҷL�@�l�[ ��w͐}J>��"�� /i� /�cI}'��
��r{�[E��<Tֶ��_F%�Al����d�)�����nw$c?\qS��l���Y�rA�]��O��з�,|����2;���_f.���� R���av�L� J����N�۱��d����c�R�P�|��VFB�3�?�mX�Z��� �k}M��uh�9Č8^��Q�6��0�֏uim@ �w'߂j׈����'�[$~>��w�[�.����d��{R�=n9TqF�����m�*�͎	��pw�����E�>ս���2��I�~:x���Ѵ���S ��|�����T����eٌ��9����&[���?-�M��W�R̥X0��px���ؚ�^�{ui�Jɼc���+��g�5-Nv� "�s�Ͻ^�O��Ir����ƹ�+���Zd�h[�pU|�8�N���GJr�� N��xf->�ˍ7I��R���׺����Sϰ�yX�OC�/fTWa�����=�������H]ci���kO�`��� 0Ϩ�\����,��~m��/^��N�ǃmmcK0ї�v�ס�
�wZƟ�]�ck�#L�1�5�w�5���A5�H3��2¬r	�=k���j�L��� 7���?Һcm�I�� �O5��kOY�@U�\�k���9�z/�-Eƣg�Rr;w�iЈ�����N�~�"�T|�y�+v�����p�lvl/�ұt���k�c�?�]\I�H�(�/N��\S��u�N'�~�E����2��x�����i�B�E*�9O��|����U�/�1LK�rsҽ��:T�y��Lm���"��Q��6�E�B�D��������ׅ#����[?yb8�ھ���b���s#
��Sʵ�~�
��6�R��T��^��џ��3IpNxq��9p ��U�o��s�i섷!^�C�vL��~]��`���:������i�ŅfU�k�� �Kh�ɏ����՞�fk(�9#n���ynmk��|m�.��!8|��������6֤�u�\j�R2ǞEz�� ��i��J��P�jE���qsJ�7	��W�,[\�|�4�7́�Ҽ��Z<4o-�
����C��!v��6�;��~w~؞���Z�<��uQ�'��+�I$6Ӓ��_^��7�4BRI��{�|���3���5��U�1,�#|ƺ� 
�2^\� ʎ@�rѯ�f_S�^����Yc8 u���i��N��q��S4ywF2����kyNi���6�<��*��N��I�sc꿅�&�S�!Rv���N�lGq1�x���Hc�'���-SD{-)�q.3�ªV�K՞=���P���*T)�>����o=rib��@#�}Q���}Ķ��	�� �c��V��(@W�#ޝ=�q�G���G�G~��v�u�U;sޙ���w�AB�6�Q���6�}�cz_�4a��ǧ�5�j�mlX�0>��X^��J�v�{��B�ҹټV�1�J�W�!�Y���sھ�]6�����_/��ڼ�߆f��b'��$�z�����28cPX�:{R��)�ƅ�-E<v�Yp�lv���|P��E���|�=zW�Y|�OC�4K�Fs�� >�W���w�g���d~���Mh~|Z�gyr�b�U-b��6@yϥI�\�/Q2�l��k.�n>�����_���߉Z�q�mǙ���� "��ּu�����*���_|-�%�m��js=Ģ0�`��J���\���oe;n�h��7go����Un�aT䦏��"x���ڛ���p�>��<7.d,[<פ���-Ƈ�=��ʹ�;g�t�|#j6�Ο�7v��)�r�绽�:k~�O��Ȱ�T�b8��}o�� B�9��t����zq\xy<Qu7�k��Q�]�����"E�H��h{��	��x�I��6�~�y9*8 �� ]|-ax Y ,�0'#�� �?*������&y��OA� ֯��c���g�ן󚬵�FN+�5�� ���?�6�ɪK*)����|�涀�&� ��{���g��j���r{���RM�r�E� �?� >[�;�;#���@f-���r}k��iᘖ;g1p���{אx��[̆6*Q��b��}N��=�����5� i��bh�F��� O�k��g��]4{�WF0G�ڸ� �:���(5��X�����{�s��F�w���Lu��튾�0��<[��o�����HP�@����|ͤ�p�M�kW����[��� 
��j]G~��#M�}N:���3�߅!�1*�fi�Q+]Xvv��O�z<6:��'1b���0s�Y�>�&��L����9�x���Z��ܳ4��� ����MՖ$�)
������wS�ļA����3ZZ4{�8��3��wezb����)l7-��t$�vv�����:�Y�7�5�T&��E��ͅ8Ϸ͊�y�7Ryk��q�9�+�S�3�J���^�w`1$c�� ~y�i>�T*�>�����zʷ�_6>:�h �m�1{�[1�A�x��%IY:�I�~�\/��E#��P��Qv��s�O�J=�gH��^ת1�͟'���W�,��p@�+H1��sA�l`�җ׽hd7z`
	c�}iN�~������ B����h>��F��l��j&i$F�{\	6�4��N�Fe�հO�"��31(����I���� \rs�S�m���4�1f'8�Ҙ�{Nz�oݐ�;T�6�9ɧ*l��$���'��=!6�W�S�ʍ��������"���;��{_Ýb��`pA��� ���5���[���6����fF�2+v�]e��h�\'��zt��1I�!��*Ϋ�5���[���V��{������q��!�f�o�>���T����`�F~�1��k��?�X���� �<�8���K6~������C�'b����*��Ĵ�ɏ�'�����X�����T)C���x���e_����W�$ѡE����sVW�����+�6�J������U�I�N�$��9����H�rHMyM�ū��-}�ҨI�j�K�P3�-C�&i�v���,�m��uiu�UAq�Lu�5�|[����_��s����|�[�1Lcr�Gj����f�;��q�w��q-��_ksȫ��<��Ұ.� �wP�_����j���s�l�Q�\R��=�>�+3�|#���Vh�pG �ßoֽ��-�Ƴ�nWΚ3�P2 �y��u��1C��o �eʠwu�3��^��g��V�Kw,����|�&��=p�f�ů�O��;$�
N�9���s:ց&�G��������Y�~?Iq$�I�X�ON¸_����?�y��K0e����)�W��J6v>��� ��q��,yo��_��n���.g�eC�������Z�ā}yz�M�� 8^	��+�5���eQnp�WԞ��}.]��c�����X��32�k��V��c �<W?st�}8���D;}23����<}����I����~���O;w�Ў�LC�m�7q׽:��Y6��=1ڝ�3�Fz�Y�7�ܞ9�t����x� JT�ٍ��9��T���饋98��!�g"�c��`zSc�s yZ�ܟ�H9������9�q@��b���@�3c H<�5c�;���Vݼ���|��F�5-�_��Q���Ϋ�,sR�ήB�GL�<��q�u9�#[VfFv�5j�Ixc�ޡ�t<���K%�*�X���@��݆��kF\RG'� �<�z�䐲����P�gss����K����9<d���09�� ����N�Lc�	''sz��*Y!m�F:����*��ӣr�ۀ w=��X�\p0{�H V��J<�i ޾�G�J��'~�6|�'��)�^A8�>mă�)w��Ͻ1�JƩ�T}���7�����Ӭ���Ju���ŗz�|��E1�g d��|���=�I��a_ZF�C�oz�T��>�����Oݽ���;�Q��ޘU�)p�1�O'� �JU���ۇZ<��0�v���T��֏,��<����J<�wp��h�
+�ÊpP[�;S|��=��Ըu��|q@�*�O�>�� ,�8+랴G	�%U�^	�T��H$�s�0+��>���z�q��]��F ���N0M:[9A�n�P2�N2OV�N�
���>a�M&��F���Xt���8�0y<��!���{Ҙ�1?{��)��Xa{�� ֫�j��O�����m���c���S��b�����ѫP�ɷq\s��Z���HS�s��2|�߯Ҙ����V�'��=�q�S� g?���J4Abf �ޛ��Ǳ���U�wP� �tX�e�rz�u�@1�%�#�4Ԅ�#�٭�f����Ci�#`��`G&��������c�]}<���机^n9a��p36�����֝����V�! <p:S���zc��
7H>��:���X9;�QM��I�b)���v��#�Q���G+[�3���iͦ��=��F�1���4�� ����9���K����)Ux$��GP~CH�b}�ۈ��LVc�5X�����z7;�G�E��f�� ��#�s҆��� �b�N�	��=j,�H��;h̖i8?CQ��#�kb;H�*9�S���R����H�����Q�W�$tM;�f\q�V�ͬqM�xQ�*B����I���W��S�n`���2++({Xv�9�@ʖ��R�ק۸�U2.@�d�ЁaRF3ո����Z"Y�LzP#��[ql� ZVe�[���-��'B��/��&�e�|�$�3�U����FQ$.AĬF+����=�j����S��L��+�KX����G�obr�t�������[�Ȱ�[�&�4�(��U���6�s_��	u+[�`���C���;�D�;���"x���]��U��J�p:���}]��úz�ETB�w1nO�5�ֿ���x��i�y��W�I����?o�ݷ�ʸ�t��a͵��� j�Xxv1��E�{����p?���{�hl����-�g�U��[��j� ��]��^�NG5���dkh� ���F:W,�:�M��m<�gX���)�S��_��N�x�����k�4M��#�=8�[�K[;Q �h��r��"�6��x���^��
��aU�mXA1�J�?�{ÿ��m�S n��-)lI��?�oky܈����_ ��O�7����7�'9��]�K��� b�|���!d�2�"�3�_�~6�m|S��y"S�G<c� �� �n�1͟��������#/�H���3${WE���j�*���o��]�H\�[h`�N7�J�����6������g����(� ��#�k��7�>�t��ߓ�u�zW����W�ge��gO��u
Xm�nkڴ=�I��8S2�s�3ֹ�؋EE���+��V#6	���]�3{���k�|��P��h����,l �5���� ��+���K����P�9�eRJ�ڌov~x��$9V�s�sS}��� ��`ܨ8�۠��������WgC��V=/�ΜuhU�<�Ծ �ZH#�\u���i��B�������E�6q�p@�^T�1�NV�ISnE��E�l,�`:�]7��&�u����n~���>����ֺ�?V�N� f����a���|%j_T���8�y�{r�1�����Y��^M�<Q�<�,s�zՎ��h���,��b�!c	�����ji�g��p����� �_ۏ.I���q_r�ݐ�~�`��*�?�M|4�c�^03]1�uz	r�O�9�W��9�����W���)�C�`�5�_
m弚4w `Pђ=����kp��j���)d�%�����{Xda�=+�4�*8� )��W1�|-𽮇��l_1�&���Ib�q���+���P�峌]<Z�֢`�<VN��MY�����|+<���Q�� ��W���m��p��I��y������>>x6+�	�02X�W�>1é��������S�X�>h�g��"� ���`ê��� ��U��)��#�-Ɠ�l��<�x�������S�� �u�1�������MKj2e�׃�(��hFH��}��_�6p�ͤ��ʦ�ͯdE���Mfq+�k��ŀ[�0�[�:[�����6�qw\�x�5�����K����ׂ~�_��n#К�G�6R�Qm�K�׋~����G�i#*Y	S���V3�S;kc�X���£�e?��\[���x���x�� pZvq�l-,���1�MtE���;�v�>�gu峈f��k��&���_-|M,k$�1����� *����4�}6躆h�)�u��+�τ?'�w�x�k��[Dr���� 
���'����R[����:}��os!^d�� �q>����H��'�8�һ�|@��ǌ�U\[Af�r@��u�-ޕ��R�DE#,~��%lq�2���g3K�7�%3�����?�T>*|3��tߵX�#�0�Gֽ�i7���[m��A�x����T�#J��n�bC�#�q�8;�����>��4�m7V���t��x���_������b9�3�~��sm�=���F��� ׯ��J����U�#�\Yd�{ltb��b� ��߱��_�Uī���8�,}s��Y��7e�gҽ��iRu��{&6�G.ZwF8e�+3�� i�_X�"���x���9��0]�c��}5n��
2���z��Y���Br�g�P�'u&wԡ}�9�a���~8���2q�+��?_��	+R0 ��e��i�8�h����,\9l�XЕ��+X���ʨ�~�=����w��.��;���_�%����t{��߶��:�0v��(���qQũUQ:�Ir�	د�I^F3��]^����$f8���4�G��m��+����A��`�[�O��sV���Üg�*��F�uT���ڪ���J�/��n��-J��S�˲�����j�F��R����.���"�X���:ʫ�O�E~���1���6�P �0+��W���vC+1(�ҽJFHWj*�W7R���i}MM��A�枭�/�H�e�H��@�.������Ic�3�QG��������O?�x��>�9�?1�{.��f����x����>�N���39��$w����튕v��Q����:7${�kK����R+w�I��:�4*�#� 4tN�5=�Q�Ҿ����a�?�쐀|� �|��k�l��p����	~-���7���Y�3�����I����MΊ6oS� �WcuD���_�&����x��d�G#���.zs��k"~��OKˉ@II�69�{���;֎�x���ų�8#��Ҹ!���ڑ���|��@xK�_�cJ��[k[w�azO�Z�}UR�G+�k鏏���~#|B�5�:X�{��Gʼ����E|��-*�Oך���h�� h���W�Jm�\�%��7^���� վ1��f��s��M��.A$V����$�_4dg��o h�7&�q�q^�_��`�� �=k�<3�e�D��#��d�r� ŭN���yv��W�g��W����' � <׼|`��������9$5?�xL��M�x'�q��Lv�Aq��Ўk��|;�"���q�4>c|� �t�^���O�b��L䁒z�J\��J䷿��3�2]M
�yg��pٶfRA�"�������Ło����|�墱�=��*#&��Qz��{�i�zt�@�[���?[��(�A�ﻍ��>��ZZ�����zW�t�]9��#�����U��ϡ��xG��l�E�)�������W�Ѐ���}9���A��&�!'�N��W�Z�"�L����E�jģȬ������C @'�=~���>�Α�,ch����}���u�F�7�R��W��>ä1+��z�ȥ)$5�{ϊ�f��s�{_�8c�������;����~px����w�Z����2�� �ON+����}rO�ze�gh������ ��|	��B�[�����L�3������*c�-�a�K,dIrI�N�Ԗz�ƞ��6��?�"�F
�銎�9�Z�Kyy5�g��= bH�ֺ ��Z��a���=?噼���=F+C�����gp'Rk@�=�?��m�Xb�渍{�sC�H���+��:�'�-��i��cv끎�sKo�B��A&�7��}*-"��k� �Y�6\�
��%�x^���vc���c�U��K�b���\���IuL�N���Z���+I�̣.���Z{����T�x�i��!
w9���aT$�n[� /֨E��3�?Q� ֥��B��c=j��r�1���q���˯4�8��q렳n(s�^��>�'� t��_�Q��#pG4���d�t�;ӻ+h/��p�[n �\�� �%�.$��˞��H��go-�ވtr��Sت�ێў����ϥF���2�@�\gvI� kˡ�_3!�d��S]$3$ܙ�jC�r�*�=��E&�,)����4� �VB66ю1�iG�Dѐ@$�.�����Ƭ.�t��5 oCḗ' ch1�ۊ�\�Վ5���v;�٨�Z����bH����:6�g��|2��;`/͍��w�)/���7��/8��S�W^CB7m�N��J�q�`�� ֭-?I�>dn�cn��)�����|ބӛP��
 v��楡�G0�e�W簩���u���Pq�� J���"��b��8�SἸ��G� dm�S@��ћ�q������$�0�v�9�8���Vc�p*�]}��]��9�i������Gz篴�->�K|��͎+����2�7,G�7���&[ށ�߶��f�:����Ү5��2F t�f�U��+��
c�+7��Q���K[��ڪ8�j�}��9���bG���b��rO�ZIO0�H�i��3�B#S���4G5���#޹S�6ߛ�0���K���8�@���F0in�zUfԭS�_��\��e ����ORA��@� �!��)��y�^�o�F��(T��9���|��]z_��!'kzצx������Ŗ��d`C�W'�@��x�OҴ�E�ae`���J��V���2D�����\Tw�K<���1��9$���맺u;�Q���a���6��,0 }��*6�mYJ����k�_��;c��H�wi��]n�nFz�A��kO�J�@>�p mJ��J3��^昏B�u]=-��A}���?&�쑃\�n;�<�sC�\��6�����q��zWП��Zŋ�{,q�������}�_+,l0��k[�MQlV�+�#�[v�n�=�zƑ�x[�WZ~��*�hJG��#>��\"��v0}+{�)yN�c�pO���\����4��s|��4����H��o� ��F�T���Lw4�R*�+��MFE�*��U=��s�)8<�4��Ԥ��r*F�]W׭PVě��8�Ҵ����@\���7!�W�kj/��v$�EẐ���r��r(rNVM��8�=i$�%^|�=FMT$;ۂz��� �P���@ J@��?���AS���)Su�0�L���1��l8��ڛ޸�q�Zhd� n����z��S4�K��ҝ$Ŕ����$�����'q����<�R���QQG���ңi.�>��u��=�!o�q�V��F�4j����]�`a�1E�Is!f<��+[�d��L�h�s.��i'�~��cڃ�3�t�Rm��O�!�iU~_�穦����IO\��>M�qޘ�3۶qH[��s`�z�4�s$.c�ʟ�M�v��O\�RBfr��=*�"�L�����jk�%�ǔ�n
q�*[u��9���y����9&_-���F9�o�5`�霁QMq(��0��7ֲY�C+��F�ӧz��dl� w������y��N㑍�b�5��3�����x�ǭH��$���w�& �Gj��d�c�i
��?٦]�_Z;���H#�׹�7����MŊ�^A5�E����9�+j�R(wǡ<S�h}����?Ҽ����Z��L�&� ��_�_/Iug�<�)m�N8|͓��|G��֡�P����^��C��1��(wm�+�t}^T���;�{g�5ϰ�g����Y�]M�}k�A�� H���%�G%����+����i�Э�U��[����W��'�5��d���c��o�x?�!�FK�}R�E�U��4ܪ 4�x.}����wzr�Z��%���ܣI������w�KN��Q���RW|nf��;K��ݵ�f�O�����h���f��z����$�Z�g����L|E�<��\���&��ݣ�-�.ǡ�����R�����2G�WԿ�8_x����y������������CP��%�<�T�9�J��:~���8Nںφ�,��{�9��_��`u��/k� �v2q֮�n-#*)s&Ϫ<��yaj�<׵xs�i�ku>��x�|����QZ���9�5�|ZҴ����h��<�����U=n�h��W���/�9X��@a�Ұt_��|�?,�y����ƍ_��"��yZ+er-�B6���q�>�� �\��|uucv��;s�'�{эUs��sX�"O�P]ۖG#�����.4Mnfl�Q���b����Z`0��^m�?�
��[(��#J�I�&h����U�W9��O�V�߀v�Ҷ��� %�>�/�zd� ��^���z��wB�]� ��9��ǅ�F��@�;���|i���t�Tn	�s_D|?��k��n�I�3���vN\����-����-4�>�j�$�����_x��C־���,������X?h�;��`����nA\�D�3_+�/��������q#n�8�|�L��:3��>9�V��̣ ��k�-�E����\}8������S,�$��{v��H[A�2����3�^�:~�$�:�����~��0MJ��%�' �`�|��Hr���D���&��M��8����8����k����I^�35��m�{?���ǨC�}�����	Ƕvz��4-�l �y�f�
v����lm�D���V3�	�k����
�^e����}+�|?����st!\���?���/���ž&1�\0��6��R?�t&ރ��n���n�����)��_K|�u������k�r-Zxn���<�ȯ�~ ~�K�ɥ����IP�� �kgmE��h}{�Kk�|9��  �C�_�lK��g;�bI?Z���e�	��F�3�G>��m[����{T�4/�$V�-Q�D��T�K��;�V���wY`x��t�{ݼn�j�Q��K]Ov�?��o�ZC�f_Ԋ�n:�@�m��K:��q�~vxW�t>���2c�Z��_���I7�M��"ڪ:}ޕ��+R�����+��Ր�o�!A��\����˄����D�g�&�v�w�K&>�)�W?w$�ϳ֟O�&l��ֱM+��~���~4ҵ}���HݢU
���V�y��O��x��0N���߁��� ��q���f�>���b��Z���e��|ʯ�I�ƭݬh��?x�}⫻��P���v�YO�M�fY�ڜ�V����Z$�v���o��\]�?��I����5�E��i�Z�ݸ㱯��_Gc&��)�������4a��;��\F���ӣZ6�>�����>�yv�M���<���@?:�>3���w�O�5��3�s)8>�Z�{���vv2i�N�QHn����o>�=���K4��ُ$�ָjU/�R���6��V]kL��{�'-� ׯG�|[oq���d�NKf�54O/QWHS�J��+㘇O��8���,Vse��=��O��k9�0!S^1_�X�ڔ�IrX��}�ѼW�$���<�S�\b�[+33����N�Q�Zjlƚ�Ew?Q^��6o�G�2y�� �pj���k�3�kkH񍾚p�U�^��Z��S*SP�Ͽ��A�A��I �ҽGR񆝤i�A���B���@��&�=�#�A.���&B� ��t��������d�읢�A�
�=3�|�rڞ����*��@�E��4��e���<q�7g��x㕦�|��,Ǌ�X]I3����t���}�݃�ɯVyu�h���z��E��g(U�$��0���j�/�,�շ�'o�q\L?/-�HD�d
W�s��Ng��pp�2�W��T�)GC�촹��d��q׊юԫc;rq����zXm�6����Xr^/��� ?J���%Z��_���I6�u�M��>�'��A|���C�6B��遊�W�	$x)��I�{�Ҿ�� �@���e�o{CD�P �1P�FX�ڋ}�a�S��rjB��#���$+��FTi��z�"P���M�b#�sI��k60H��@���R7��wR?J��p�,s�ֽ�Rm�m�'��^/$L��N����L���Fz���<��ZB�h#�� JI����6�ߒ�}���R}�$�w�)����m����[���)��� e��ۜ���:�6����T��{�<;�ԯ F�5�?ŏ��o�g?����ݴ�/���Y���
�++��|����Rլa��VG���67ڔ�b��g$r�I��]/OKͫ Wѿ�_���[Cuh'0�<��"�R�WY�_j�{��I�㚨nFi,�������+����M��|E-͝�F�G���1� � :���~����
�ϙ\L��o0�����a����q��@�; y���7�5|�wk#}��k�4� C��+ ?�������Kcp�kKX�Dz.�-����'�[m.W�����&��>R) �H����_��3V$�ZFVaǿZ�yp.��,���u�S�<��>�G����R23�W+�� ���'vp�Ozܼ�i
��.v�x�k9k�Q�v_<Y�<5���!��'�I\��w���u$+9 ����5mi�-~�Fe���\�������l�{�4���>?v_ӵ{O��q��jF�L��������#�~i��]�y�N� �+�����)m�ߥeRKb�}�O���|A��.�6$F�p6�2}��u�Z�	'�z0��9���y72ڗ2��������[�,�q�ڵQ�!��Mf��������mt}<Eq�m �����|K���)rr;?�z��+�2���qYL��s������_R��M�����q��#�#���0�����8ֽ�R�hm���ȒQ�?��x�4��uD��L���UL���^��wu#ۚ��U�����j����<�¶$L��8�ex� ���
U�=~��2��ڀPX��3Mf�22p	 ����l����d�P�v$'8�� ���� y��,F8�8�*ƪ2�I�Ҁs����99��`��i�śoM�?� >��ܑM���Gzn��\c=;q�{�0�2pFO�L	a��,�q�CP��(�J�Pz����1����I8$q�<����� �C��[���ە����\�ǽ;��F�s�қ���Z~�۱�i�v�����	�(%G�*F\�'��M�\ >\q����y�"���n�zsK���8Α1�$��杵v�`v�0O�I�=�Q8c�^�QC.
O���(X�Q���(��Z��0q��)���Xә�N9���6O֔���'��@����O�P{�u��G��i` ��#�>�M ��#ifO�x�d��8�)��ON*6!�h6�S��RC����L���zԑ�v�n�Pc?�-�=}�&r@�n>i�>�����1Lc�!�<b���pp^i���>H�pÏ��ڐ<�=��N���H9����e_�ՏSҚ�|�a��<�� e���J�����zs֑�^�g���>ޔ�aH�t���i���OϜh�6���6߯�;i� xQ"�m�r�Үy�T�Q���iwH�����J���L�W�8�n���E㚽�i�M�>pw�v�q��߅ ˑ�zqJ����c�3�@�
���#�OS��x���{��lCS ʰ<�$Rm�u�=jFR[� ��>�����^}h=�ґ�v�I�8�33`OZ{*��;n��j�p'��d�A��K�����q�f���䌌sI�h��{g�9횉T���� �A=;ޓv޽A�IA�?�4����M0�p��AI��-�u����� W���@
�2��}iv�.��k)l��S�� >� �����d�������T̥xڤ��I��D�'9��1w0W��zR���[���P!9m�b��>^=��� �R�ށ��Y�9�=�Ѵ�Hb3���r��8�3�HDk��t�I,�g�֝�v�g0�~��灊�f��'*�t �������N0GJ���u��_��H��d9�AV|�̹�^�UU�v����VUJc��L��B%��{���E�֪�#
�FB穥~���H�@I�p���TL�\g�֦��^G���T>f��R*�cx��fN b���=����P��Ræx�fe\���]�Г�T,݀��O�?Aӷ5{M�LSo�ߜVv>^��Mۆ;����x�m���=Ko� �6�lこ��^}5����;�4��|� P��ƥc�&��x��r�Vpk���&i�Wv,ܞ:�L�-7g����O}��zR�NM�C�A~�Zױ�ĖQ.�q�\�\���5�������CI�0RkS����nF�flq��-�0[�}3\���"�XdqP����l�e�n_��jx<d#����m�yv�
��B�E!�J�Q]����k�=s�a�4�k����B�ұT
I��\�#�z�y����S�[>�>�;�_��r�x�FR�I����N�ӯnx���~���B�7#��in�su6!��Ï5� ��3dg'ןƩ6�����SƎ� ��K��s2V�[��I��"�����qӟ�Q��0V�ip���>Q]�� �]sJ�ҧ��&�n��vCT$�Fl�Ҕi(����I�KtR�������R`e��u�7׮�j�i���M�a�\SJ��NM�U�ėq�6�Zo_H�,��N[��4��ĩ����\�\�b�����+x��z՘lBr0:b��#�;y\�� :��a��<�Cx����w�*ս�kd���6c؊-q�2���TEڳH�#>�A�K٘��r{��m}�:u����v�t���f�9漺�NN���׊ۃ2cӊ��c�L��5]��ǥ2U̹5��r�OԜ�#����e'ڵd�'`T`�v3�<Qb�鮯!�}qQǪj
�@l�s�k�����V����D',��u��[R���i�o�֤eB��ә��LWg>���s�ߝ*Yܷ��G�5�$��҆ˮv�=��dr]���ҵ����a��ZH��H�7�l�9�F���G�%��K�
�,) ���B�`T[��0+2���G�N��� �����n��Jw=q��������-�a*��Ү��K���☊dY�9�Ne�2y�Wv��3�jSf� E
Q���<z�� fa���t4�&�� �}���1@j'�GR?#N���W�9朎ϏNƜ�>�#��@��M-���ӭخ[q$��W�����^w��m��K�~CŴ}f��) ��&ӏ�d�70֦�O/��i��M�G$��;��4{��F���H��Wc�c�'ֶ�g��Է56W�w"�d�K�!�Y�06rX�ʯ���ϽS�����?*��ďп�.4�����<��1�־օ�Bu�|[� (>e|�N��+��[x����n·�,xZG/�45���~�+ �o1���#a�j�l��ԭf�h��6��q�U��mCc�3�Wo���WW� �B?�\��q�h5�[^i�`������5캆dӦ�yܢե�W�9?�5��2�r��~R�|���#�P�i�cZ��k���֥�fi�I⡍�JFx���,��_c�PI�x�t����R���~)�`�<C�:�����tb8����߅|�tۜ��� qW!��}��3�������W5lo�y��8?�}5�4�D����+�B�m��o'#�~5�x]��>o�MIo��kyv� ��ED�Vaf}s�\�r��#x��-&H��H���rs��Ҿ3���ES��\V����9�N���$�KY$\:��c���^h� xq��jtp�d6x>�0�|��G��ڊ�5�8�U�5�=�94�A;H�?���x��W:����唏�x�k4�Ǹ���� �O$��r�r��o2�)�ڙg���+�m ݴ���M�NI�EL�z
Z
Ɨ��]w�ۘՙW;qK�x����]Xv�d�ky�Y6�8�k6���_�O�+F�����pzW��97�s�WG�$��.A��R��?(B1�ޝ�%�x��E�M��X��~u����,'�%�E+����J�Lm��I_�)��ˌv8��R�ܵt�9���I��m�.��ƙ%������խ�+��q�S�ڬ^���>d.Q>����j�0��W���ۘ����Ԏ�����:G�;���]g�t�[���|�^g��{sޡ�,z�#�� ���.�����I�����Z���+��c`g��.2K�+{V���Z�bM�n7u5O����oȥ��Z��9��y%���⧎�+���@�y�nQ��i0�9� f�\�l��4�̼�Ա�u=��5����U�3L
C,ʣ}E&iی�7CD�v�[>�����޽�v_A�4��[���RJ����Oަ�c\�h�v�8��Q��'���Hf�nVh��c�wz/��x��7�ӷ	9]Ǔ�M����zqMln�75�x���<qo�c$o�x���+�>�<0��]�<pL�#��s�� g���ɨ�l�%��{����}sZ�d���y��9���g¿u� o6V�&� �Rzzz�k�C��T�ۜ`g��<��Ev�����r]�Z��9 �����gIP�!��޴X"�J��;ONi�,�9��֗��#�x��+m.�[�n��w7߳�4�3pt���.�}r����ǚ2�W@K8�K�� ���������eun�]� ��+�����Z�����C܌�ʕ���Ee�A�)UV5�q�i�����X̦9ն�'�z?�g����o,�Ym�8�C�;PM�8�����:zR����a޻|�?��^�P�f�KD�����\4+%�,q�\��<�@�.{�J��\�� i����u��v���b�ud���\�7�g׌�X��EU�!��M�Я#��M&�m��秩�|U��Y��s�o2�+�#4���@R��y^�3.v��2+���{�Z5֧e�� �c��=��*��_�~!��qu�fB�d�}Nh���8����=�� 潞o�'���U�F���ߵyΟ�� Z���b��K�}��~l}(�2��f����/�������Hc,��>�>�潳Q���gt�ImFߓ�9�yG����T6:�lc����+���F���ӤX��®i:T�ƭ��fY�8\��z��K�n�j��Ku`ݹ4�lM�x�Ф`�h����\W_�����H_P�yS>ԑ��]�g�o��u'TF`��q�l����atyW��OoJ��M���x�|����Y����T۱�q��� �!��i�K���v�4r����3���E���/x�����`�c��^�~��)��g���D?�YA9�J�; k?��9=�E��U) 9�=8�阅��;x����v���k��c?�s,q��U��}1�yGď����}Ymu%;%� V����������.~v�8?N)�7��RH��'����8վ$j��M��//�q�$�����j䎿ʤ�FRYin��a���Ex�d�zn�}k�վ��C���4L�c�B=q�� ];̏:�InX���{�i���~��������?ǥj���@��o� Un������/麬�d��B�䑞�R���@G=�P�r��G�^����W\�N�o���p����<Z����8�����&�!��!l�w���̶<�c����b��X��!f��A����� f�{�%��A�@8�� �8�F�Q��u`���\Q�`�W�*��u�K���u��R��>�׃�hz���&;R���6\g8���R�C�V�H��#���R�1fV�G^��9�W�?e� �~�W�+���]�q��Z��/T�ƽ�kk������`RL�]��oQIC�z��E?b�JH��*�#	?�����O�����"�au8�Ę�2v8���4ӳ�޶|�[�x�*�&{�[ v�5�Û��|�̚0�(8��6*��,��?��K}�)UB�`pG�R��\0$t�[� �y�\]:���0 ���Ð ?�QɄ=z9���^��_�΍q�1�B��<g�5����.���Yj��+tʈN��W+�<�9��i��� ������j��� ����xv�R��[?9w��<u���T>8�����V��"��V�ǹʦ>\g=yr�9��M ��N�C#�J�� W�� ��5?��2^[{Eb�c���k���o�iS\��+<JX�A���{S��9��|��O RK(������Sg���K<���
~
�?.��Z��I"�{*,6�U��E��4�4~X�s�_H�_����I<W0��Kd��1^g�YO���>T�_(��N�;}iىI5s�󂐣�Tfx��_MC��5���aIgj�?��^s�c��~�^�~��d�q���ÙO#0I��j/0r;Z��~�z߉4�5	�Ȳ"��=��k7�O����Em@�,�Ǎ�/\��Q�Ù=#V
�r� �zt��(#�^k�>|��%B�0.�x�c�8�g�vڗ졨i��$��Z���SO���c��#-�����~񰢖��m7S��\	avV�<���
��{�$r����M�D� � ��K�\I���I3Q�H��0 �?���Tg9��S�'�����֐yl�T�sϽ7��Yx�Oz{:��jF^ǭ!���c<qQ��-�}�Rc�QJ��q�ǥ 'R; 9�Ok��g��*���=3V-x��9#�>��Df%P ��LY��@����$c�kHثD��o�� }S��T���U��`v��QyȌ#>����d��:{Ӽ�$x(�z摥Fn���Z�n�
��z `��������?!S�L�9?�3T�� 1��g�{�@�����sR��ƣ�֫r�p_���R��s1w�8���sN�5��ޙ�mnO�F���r3�M��WqO�2y��׽�#�X�����aLk�Y�j�u}�6n��ZY	�3NV�
�x�$u��FG� ;n�>�Jz���Dy�43�=�dV8�U�����0P���=d-ߞ�4�#[���/�*O8���&�6qU���(@�K��ɦH��~��yķ9�U���=} �/�YXv�'�z�>k�[�Z�E@rp=��?ƛÞD$�ď�G��;u�!�m�2*x�V�n�Mdػ��j�ƭ�HBO�E��p�\��x��Ǹ���-n%��n8�s�j4{F�r;P!�C.{S�
������.rz�v��1.���@(F�4���rH��Jwrv��Oگ��&����#�J��F߻�5]mæ��(�� *�vL, <���hKz��\zQo�#ݐI=�����%�c���ř�#i������_��6��O?Z`bc�b�s@��v����pi�Ʌ�dv�U㹋`20���_�b�3�Ch'�d2[����Y��޲M��ws��!���8דϯj��.�`�!N+
k�\�n5����ǩϱ4��a�g=��2^GQSH8>�`��;|��۵W�Wq��8�Fe��+6K�73LV-����i�֑��I�85V�Z��e+��g�w�f�$���c�k�)r==k>MVI� �O�f�t���;�l�qs�c���;��LQ�<�z֌�(Iϭe�5�l�z{V�$Bpx��@�PoD��ɬ؈��� Z���%���ڮ� v�d�Rw?B?`<����F�?���k�}�hS>��_��!q��S��c�8����$A)��-���#�0'�(�Қ�@3�R��Ekx�M��
�3|�~�����_��_�4�277�[��h ��T-���&q�?J,I��t��6q׃���ogi#��{m�ll� 	���N��>Nܱ=}�V��&E�d`g��+�� �J�w�O�hLEhd&O�1�R.F��t�[��0:��o֐���[m^��,1_�_	~��x�e���l��q��ο9�3∴B3��'"���O�m����c;���)u�1��T�icH��ɩxFKh�#خS���/�?�%��֤ȱ�Hs������� m��v�r�S� /�+��?k�[H��]���`J�3��N��6���muۥ�< f�� 
�h�qt�p�I?�j�h�Iy}y2���哃�j�۫ż�n|��v���i�F���WE?h���tV'�9,"����8�5���̧aޮ�'�#.�pF:��*k�G��9�U�Kg�v5sI�˫A��^�g�ҥ�4w�iv�̶��s�j���kXu{�۟*3!�L��bү#Qy���{�T>��Z[ˉ��$F�L�+��+�R{�}'R� �������6n�=�FA�kI�n4�Y�1�y�y��]�m^y"��3y*���G�.�W����5�!y?ƴ|M�H��%��2�����߅��kwpTU�����*_]�v�L��-�V��s���W�I ���p�ۗD"�����j����O���9#3�6�*�������R�\���l	��9�T�v�X��G0Ğ����ga򣓓T�`�!70��º{�[-cK��Cǐ�x�H�xu%�����7`��?�Z6���"`U�2Y���*��Ac�<?mڑ�H��\��v0�oi⇎�đ�s���d��+�-�[YQ�w@<�����2���� r0H�Y���l��. K>wq�0?U~'cϰ`�
���<��r3� 	Oά�����F#�1c����'��Қ$�m���~�甬����%�2~lR2�m�뚠f+!#��ʦ����?*���=*2�ӧnQ��t��g�R���
n�x�Ү�^�����žU������iG u�%\���@��0�6:獬"�O0<���$� J�7��U�[�J�l--���F��䌓�N��z���?��>6�i[o��b�n1�ע�{�E�x��厥aj�aUw(�A$�} "�[\���_��<E��G�h�̻�H��r�� LU���	-�S���A:F�"����~�ߏ���W�ĞEY��
69%>b9�����rxo��(.
!���J����Ж���v�W��z+�l4K*n<1�E���A��/K���E>��ډ�$���������F+��-ޙ�|��ҘF��J@��sǰ'�x� �}S]���X����Qw�$��ӵ�W���9�׏Χ�kv��*D�&̎���?�|I�M��➷g��;������;�YkZ߈5��$�z`v�.��~�� �Ku��m�����^��fʉ���I�����[t�핀,���9��W> |~��c�ˋ-{I�=5�,[x,2Fs��w���K���o7��= ���|[��t�R@l�kf!&q�1��S���_M�������h/��{�C�����g�\�_L��⇃>�k�y-�{�T�F��\�ڼ���b�c�j�Di�m�]����c�*����P�'�d���@۟�V���3�>0|$��R��d
�h�)p�'$~u�~ ��;�K�<9�����YUX���v==k������SH��V���3=C|���߅v>-��� �6�x^wy�D�4�l�'۠��L|Ϝ>$~��x����M���������_6�.��Ic���PW� -^��ʺ���{�k��v��l�����=?:���f��O�I�����T��ti%����߆w�&�#g��ᮼ� #P���|]���ׂZ���4-3�À3��_c_�>
�F�'�l��=�嘌?�|)�P|m��o�!��?{ecq� ?37N8�֟��-�  ��:��6:��o3Ƹ8�u�Oj����]����M�m�n �ι ����9�'�����.;fS*3�8P0zsҾ��[�r��6�-*���9��OG�/�j`|	�o7���+{n<�b�~蕪� Z��|E��O�[��rFO >����}�{���� �zĒ\ �KvTRG,P�?:�?gֵ�g�}kB��~�r&X��"�~h����o���Aj�]q�jJ�?޶�q��}*��.4�'���O�#��	���Vl@�8�U�����񆣨_�He�=�[;FG�+���2�(��|D"�kY���E8��������<�g���t�H�I�V �Xz�:� �����Ɨ�(��-퉲&�c��G#�־��ޓ�]/Ű�j!o4�������\�� :��������Kh���P��q�u�~U;��ci{�kKAJ�26��o������Ox�Z]��l�Y5�3�\�b�=:q_ �-���|_c=��q�"^s���_�}��S���w�RK2�b���Ʃ-.�=ϝ�h�c��</�Mw�}��M������8�]��[⟃��Pӯ��Y6�S��Bx��]�q}k�|*��M�{9��F�G����_�F�⟇'�֩���%q�m+�(���&}�*�g�~,iz�z��$�аܠ��1�z~U�"�;�#�QCk�i/�10!���9�u��O��������#v2H8���_��>*|Y���ۤKɌeO'/��� <�fF��������8�����q�_\��X 9$��x��Y^$���/�b�M~"�;�E�0�w�!H���?��'�Q��m�I5���Xړ$Lރ<u�&���Zg�jAo�,v��ۗ���� *ad��� �]7��|9�˥�
�����\�+�ګ����<Eck���g%���y<g�W��+�o��ۛ� �hyWaQ�{�+�m�t���0Z�?�Rl|�<g#uL��������#��nk����-7����#A�׃Ԟ�����7�!����v5�/�1�->��X���c��U��� ��T֚����|G�EM��)�5���G�s�W���8� �<'�|����+��{�2�/�'�VD:K^��K�x%�`�s��2+��%���Wx]Y��}z��+]2��d���m<]�{an���:��Q���_��;?�~��/.�̃x#X�z}N*׏�4��w����n��7dd�� �.���״�S�~�$*��Fq�s���T%���t�./�����vX�䷷��n
1��n���7ď��>�y�F^kTh��0���Pk^�<e���C���pZ9��۟�+@h�|'���m>��#{$/3�V�=��j~ui�"�"��%�ۑ��J�E�Y��Ɛ�M���2�� d�?�������J&��� ��O>��߂���F��j�`���t��6�џ4��������KD��/�Rz�~bt���4�sK�<e��e��� B����?�6MJWľ3�Yngfe����rI�� 8���o�,t� �>(�YT?�0L6��F~��4���^����w�a�k�Z��m-#��#�Gn���z��?Y|?��.l���@Qј�d��������ҳ~輡rq�'?�{���]'M��-�us5��l��e+�Zj̖�v5?h�s�~�Mf��ɱL�#8 �pGz��gƫߋW{L�V�\g,{�>��>4�;վ4x�N���[�I��
�K���# �k�_ړ�^����O��J��Ni�9��)lkN�-���7�,��0`�P?��ȯx���f�ϊ4�ԣm���A���<��?���?-C�<�D�=��?_q�j����=����<R�"~�5#%��?J]$ԏ��%�,����V�,=�}�}C���6�y�Mh�w�<���w#5�&��W���w�����B�Y8�����5o�V7Z�X�~l����N2�z�Ư��x�➟��U�1&�9�8���_�kM����l���}��:�� �z6��Xx�3P[���+#1�g޾r���7i��|;��L�q鷂[��6���ߏ��^�QM�v��mO�o��'��nֳ�F��N�B G������\���O��]H)2Y����w�G������-{������%e�����x>~���uq:Xͷ��d�΁�[C���=:� ���zd�����v$�����5��xg���ɿڌ3�~;��׹�[�|���x1.��B[+�ΥT� ���n�s����EpJ�$Wܮ �K�=�?0��'�K��$�0)� 9�k�پ��?._NH��� Ub����+��C�ZK`����`8##��ξ����S�c9��-9�5�w6��k�~&��ouE�x��%�_(<`���5�|;�e��������G��6���}Wl��+�UW#����O����%�͛�\.�L��~����[�����x����[�Ae��a�m�:��������N��O���_�'9���O�u�1���_*�	A�<�$�}k���o>��8P�B�poO�?�;���-�<"�����}6��L(����۱��</�?į�����̸6�a��HRGA�����U��E�	�g�ޘ�Q �ӕ�s�+ش���+�3seyq����*s�u>��W�����:/��6���d����SX#�񞇥j^\k�4��2oE9'>�����7Z5�Ɠzc�3���B�1���W��GI��t���Iz%�)������:�������w\�ߙ�#��'��ң�2.z���|P�����&��a3�U^��+�c��9Z��{�$�7ڣ�u�Vݒy�nf|�ȧ��1��� 
����dg�b�Eڭ�=��0�Fʸ :S��K�!2~��A!,���C7�2x�$�H+��֍�Eێ�ϿzV6F߻����u�;b1�~n��_v\���c<�aR¿�ʜ�ңz���zS�X���A������t�R����*�1��'#ۚ�o�9�;f��K��hO�Ë�[�bw�Lv�{T`�:�5��x�M7O�b}���Ϸzd����yr96) `�q�U!�6r�O|��5婑>A�����!e@� zRlk̵}pOʤ��c��-�ZQ�� d���G%{�����+�0r~�{�g֥6�E�m�s�t��5��Ny�YR	8$��L�p�3��?:�cܱ��ii3�v�L�|�zf�Ǘ���;�ˉ"��� �q��A�8�8<UMQd�|1��*�و�.��z�����m���b����´�'�?�E��N�-��$g��o�@p)|��nT��H����P�6�b��r�q�Mm�ڠ�q�qL
]�����:��y�֒�0��=*8��i-���i���L)�j�1f�٩�5S��^E;�3R֟�)� U�c돥T�՚� v�e��뚱To3��O(ܸ��WYLr�*Ġ��1	�1��2yg�檶�4yr=qN��FmǾy<֥����
ǽ!GRi"۷��g�<�8�J�/����b����L� {�cE�5��T��r:���)��5��)�Gu��:p�☈�v�Z�n�� ��#>ܞ�%���IP�4��p�����k{���m��Zw�� ��ҥ��+{^n�c@#?vq����ҫ���\V߈5�{� [5�G&��yߚ���k1I=s[�|`@��\�%�x��]��\�� -����Uul0a׸�����#<c�}i��fg�Q�^FN3�k/��c
���>�V�����=+����zr}�5������'  M@���ʰ6� 繭[�]\@�cn�Ʌ�1-֥�D�D�@���?�lh0�q��z��D��޿�k[äI!S�=� J#�����c���١�R�g�Re� t���a��y_ư�;��wȮ�5-c�Q���$W7q���F�==��xg��\��y;��2k��6ZT�0�.+Rk��} D��^���X0C�@�w�����:�l���K#��y��Z}�g	���[�s�7�@zdq�-�+���ڬ¡�A��*�m>���V#ڬ�お`ҬQ����Y�����2dҵu�Ė�[�+"ٌ���jC��~�� �=A���&r������5���	�������>�e�E�Q�?���d��rKs���G������A�?C	A�F~^�H����}���:u��a�U��W��.�B�:Sb��`�ۀY��h�����
��6�J���ğ�8�Q�YW��k���Y<��eݞW���CX��֮L��p>��kLR܁��$�t���i�'M�8�o@���z��c@b��Jщm�F��G'���:�1H.,�y@P}G���;T�%H��s��5��=5]QQ�*x�}�� 	�B���#oFu��e)��#XŽO�����]��}���x����@H�9 W�]�B$AG�?�Eo�kh���0q�F�ҳu|���_������e_?�+��jȹ�}[�FM�7��37J�(��5�l�����z֜���2э9Yh �Һm=��T���N�̫32� �u�|g-�Y%�T�$��՛{���G'/={�[�:v�����~��(^�q��I�x��mbE�Tl'���i��+h20h��s��dz~��L�u�W;�G�����%X��$(�jOB��5�=�2 P��'9�P׮o|Ap�RDX�U��T��9/mՔ�f �X�,��m.��5j;(���Mn,�2��6���.��H�YGE�E-��NzWK�K+�][SeC�D]6� $� Oβ|[ec�x<�=������9�����n�!��P��8�r�k�Ge�Q�\�o3����l:�W$ʣݏj�o��x��zb��I��Π�n9���rW�>�d׾���8���Ś����<%��n�g� �������h�+�.�V[�睧������&�����'	"���v=+5%{X�Wm��&Ku�<p9��<'�A^��L�\�� �k>�&ߙ�#<��mxN��x�F>�ֺ�c�֤a�RWn�~`q���Q�H�jZ;�n Q��aWuvx��� W���W��E��rTmǵ08�eT���9���?SIn� `>���N��2*�@8�4��)���)}1��C��߭ 6X����*��ۈ���5Z5�s��,�<�Rz��[�✬��ҙ���x��Bs�������|O{�}R+�Ih=?�'C�����8�ӡYc��_3"���qL�:��>��Қ��{oŏڋ]��6���=�2n��[$d�Z���T�|r�K{4�-��ya�>���y*���0��px�HB�6�=�3G3�m�:k���Д�P����t�W�|x�~�X��0�h����]��B�QǧQJʌ���B�Bk�s߼]�bkzޛ-���z~�A}ſ.+����&����3ofn���9�XW� ݞ9�*�a����˘�i��⦥��TI��q�vg��^Ѭ~ں�����_f��sտ�|�
��\���5�N	��9�����I�Ӯ���mrI�4��ӅӧJ�|I��x�Mb�����B���5���`iU�@�����׉>.kzׇ�4#)[8
�^�*���}�Pk~�c��\�w�eG�Mx�m�|� 1��,�X#w�W3%��=s��=��:<�A�m���}�	8�}+ǭD��$O���-S;G�Ҕ��際���ީ�ķ��H�KA&���q�W�/�q'�+4��,?�K���ϭ;sm�4���� �O����ǀ�K7m�F��sY�})B���`:o��uψSF����@�����և�?���Y����#�r:W�|����)��*�y�wp�>����<A�V���b�d`g#�������2��?��3K�;7=O5�66�>��+&C�J|�yo��mn#��Y]��?��y�|M���X�V��k��8Fa��+5a�����cf��4��M�ZIG���c����ۗ���-��!���G��2=����3I�m-��j��<�r\�4s=�C�>&�l��(�Vד��ѲcV��t��	cU�0w.:�ʣE�#���	{�J[��	�KU�n�)����8\�y�?SG�>+k^�Eƽk/�{q+M*䰑��z���^@\�i�hۜ矘�ޚ��:���]WMkP�la�`��#�~�6�$�]rmY��K֛�2��1�&��k���}1���(�`{L��'�MK�#��d\��q�"�5[ο����嗆s�z�'��-��ʞ��ݯ��G�(݊ >��
.�h%���d{�@�
8=8���/��-֙$����p� ?����o�dY#1�c�W��o|}d�б��9IpF}�$�#��� l������.[���yƥ�ĺǍ�W�������]b�;�A�/�q���
�Yv�d`q��W3_�|M��Z�j�7��BH�9�<ַ��"k~.�m,/��K{u n ��y����I��NO��Mʹ���<I�}-t�Y�h�$t�z���1x��M��A�%G�W�N��_�)�ʸn�sU�-��Wt`n����>�k�~��IC��$��t��9�"����N2z�$��ў���[�>,�kE�h��v2���^k���y�hzl�vW2��D���kHO�Ё����)VNI_��Q�~��i�1Y�;�C����.�q`�߭:���߈?�L�oU�nc��ҳ#|(��*�wQ�� s�)]���o�E�#-�� O\}x� �כx������V��.������?p��z���'��I�cП���;�b·�]�R����%��s���)�f��9��Q�y�m�G�+!�8a�v���c���?1�n731��B����L\H�ݼ�{T���܏n)�� ��#�t�����bn98��\���.n�<�Ig���V�#d�ǯzx�\�M�h���<U�hVk��� ����Sx����y��&��W8e�ǧ���	!E��{�PnV�� P�#���-c�,�c?���+���ֺ?�?�W�<m��1'hmq� u��rG�������e��*�>_�O��ȍU� Wn:k��{�b��e�Aڣ ��`s��F��^i)4�k��q�Lj3G!V+#g"�s^���Q�K�^Hd�C����V�4�y��:m�r!��ܷ)�J��G\��fV��A��և�> �^#��,.n���� ��8�`q��t��� R�H�����	�-��y��~�q(��+�1ؑϷ���g�x㶷�"��Vkh���Ga��ڛ�;㞻��=7�ad�%�7�~��sƳ7Ȅ�q�J#6R� ��Z#��?�G��a��C�Q��zu���ߴ�<Ynl��6��0��u�ה�L�!*>^��]�������BM�L@(8�nrG^�Z�wn���&bYz�p?Njk^M1\�6N�Z�,��B�������NpO*����{�`dg�J����=ǚ��^}�����Za�֘����^N6}�1T*�s�OBE)W$�@�~p*��v� ����ڪȥ�oi�N;�4��X68�C ��>����/�cҐΆ�j� ���5b�~ny��-���Î��[��c� �VI�/ {
���ʤg+��� �ZW߻��1X7qǽ7���g�m&�T��"A9a�� ��=oOM&�Xo ���^��]h�y���_ze���L���K��4\eYr\�|��{b�4�ˑ�`��Eg�-�1��^��`��B������X�A��j�F��/���@��z��'BxU��N6��%���kR �ǎ2���#s�� &� �T�s���Cq���8�9����a�5#t�J��=p:QjY����=�)ppq�OZ�OṚo�Hf�)��=zS$M���Q�F	v�f270��&���|�N�_QfR	�*��n�:��ե��7�� d܌�:T;�\ǷZ��i	�߯4y8l0��j��3n俱�#(�qӏN*F��A���H񓷏��3[KoNG~1V������÷�8�Rj��H"�D+�ʬ�BV��$`g#��0]y�O��e��~���cy���j��N1�P�f�L@�����R���.�GP�r<�)#y����E\��_/��v�J��>f��ކ$�4�"���zv5����7q��
�ܙ�\�恑ݑ��Tѡ1�*�s8�*�2n����}��8��=+<����kKPG�A�N1Ȫ�ٲn$���P+�dEl)�x�>v��j�t�\��.sDz{H��i蠭���;�����#�e.������Ւ�cP{u"�eճE�w��3��Z�l'*2�NN[�¯�n���LR,(����:zS5hDq��~Y>bW�WM����\��:VW�@m��)���FX :�HW�`n{��[�%Up2�Tq�2\G�!]Cb�+�M�[^�o'Ϟ9f��q�ִ!���Mʭ��#�;�^Hd�<c�ᚂQ���ӭO,+������\@m�A�.qLHײ�>�I;F:�'�#��@��ҺdɈG� �y�=/�
U���M�Ƿ�q
�S�Tko*��rG^k����q�f��G�?��du���$R����Fܲ��}m�3&0rһ-�(3W>ĻB���N���������8㨭�x=|7tOnա������(Q�4|@���X��w��u8-ro2�1�{�5�6���@5�����<̎1ҳm���#p5%G�G�_��n���hc�
�N97*����	�&�^�� ���1� ֯���/�%���e�֪� N�*��b��ƬY��$H��EZ��Ul�Bҏ7h�,�s��,��)Z>��)�������e��N�k�u�#�`��f>�k�-��</C�l�^�H��V�.Zw�##�V�ЙnT���-�ݪwCO
Y�9��S�\`~U�"q�#�� �>=�aq�DW#��9jEe��ҠG�|-1��n�����ht}u
`�~���&ĶD����_mk�$�#f�d�ǿ�g(���;��Oi����z8v�M��˄��b�6�[ƛ�ݜϽoM;G��³{|��@LWQ�$��F�rz��i����c��� �@���#�pFGQ�:�eVeV�G�]-�i�,?4�ϭt�x��1ҹ_�l���v:| ƛ�=8�L��J��v�
I����1�GZ�$ar����%�F񌺜⓵������ �0��H#��Yڝݗ�n#����J�����l|�I67Q�Lw�3xf.�K�4�Y~lb�o���Vka�Z���q����W*%��P���n'���/���Sq(h�I@���>!������ܰ��5N-�r��c����I<�yj:�'�@+��t�4���*�B���@~�s��u���2�r��X���Qsu#ZN
�S��:�QԷ+�ch|��%Fz��`�J�^�=�0�Ȅp@nO�?J�)l���4lq�v��.���E��N>�=�� u5ؘhz�V����|�#��_0� �g���Sjׂ� M���<{�s�ܚ�h�[�j� [�Y��b�n���g�^0���C�4 �q���`�������2�v��1'�0O�]��O�p�@���
��������I��#=����浩��Ų���s�k3��e����� c�oδ�Q��I�bB�����2�H^	��m^����Ʃ�\F��v�2��1צ9��a��"��o�P:`�L�1��r��q���J��?�7�G�0��T�U��i��S�B�wn��O� Z�_=?�>�M�a@=:���d�i�9��iU��*3�y���BrsҀ�z�T����z�L~`	�J��n
�:�Ƙ�w`��<��8n��3�7ަ�\c&���+B����ކS�rr����q@�s����n�֝k��*B���TWKc����TȬ���T9$Z�)ls(���<�֐�|�z��[��k�ռ}��,���ITLr�$cn�s�S��j&���9���3#g=FG�R�}pr}����\���wtFT9���*�n�{q�F���ӊ��uV�B̾�V�O��lKgߚc�!���~��܏_CB�����'j7��Ta��<�c!����=8昆n;����><���S��W�ї������C����"*Fjn�����>����88��㑐�,N9,��ˏ��1�C����6���Y�ˌg�kJ	]�D�*�\�F�p1�nQ��9��M�������Bo��+�3�h�����ׁ��������ʋ3���R�z峜�u�9����NU������n�n��]���G23v�8�jE;W��5�#�nOJ���=�HO�MD�6��59��r8� ��Fʮ��#�y�q��^���"�."�X����ּ���zu� ��ٟĉ�^]y�U�c=I��U|���ml����jר�ʄ�]�l�צp~�⟴/������p�i7L����W)���5���p�I��-�$Q�����|A���յ�J���..ds������sӟ4��M�)�Ȑy`�1�݇�w�~Ԋ��00�ozR��=�u�����sJ����Un��OJ8#���㌖���hL+��jr�$zc�S�c.��a��9�8��K|�F.NȮg�B�#��=*E�p�#�a]�~��
�M�C�ksR�C�q�l��OE`룯겵���7�g�����~�8Ȯ��n��ؗ~:�W��%v����RW9�M�ѓ�Ǡ��������CL�wpNT���O�H�*�#.��sRmm�q���Kd(�D�n<z�޷���B���C����P����?�=��Ss��r+_S�b�%����+2����#�;�U&��qkq$���6UNq�JӺk;uD~p@�|v�4d�3TI�Ј��y�M*�|8�3��x�F�H��y�[O��Z"#qҳ�E(�e*�\��Fa��ֺ;���*Xd��7}�_X�2F� ����`b]��'����U�VC��O�&w�'���z��ޟ��Am+�[�|�٪�&J�[���椒�p;Nqҽ�����lLn>�G׎��� �y�l�����%�9#����eO ����&�߆���ykp�3�\�	�UrU��������*�/�#4s����@����_���cȷb7K����m�3aX����q�����v�`�G�ϭP�4��ˡ�Z��S6�>��s����uĞ{�=��jIn�O���~͹PA�FB��H����Ɯ� :P>ozp��n���Mڙ sG��(�O�@�"|��R1�p�*q҆;O4 ��?Z8�<)ǥ7�}�>������Jr�$�z�@�n�?ZNA&���h#��Dy������nbzz⚑0n$�Js��ib��`�2On� Z ݳ� :�v�Oc�o#�OѤ�;�튱o��h͞}�hF�7�,���Taә��5ؿ�r���Nj�zI�x�@#�](��1�҉�֏�W벇B/�ۭ#h�>6���94������S�p��k`�0�����P�p;�����g�h�\Ŋݥ�ٿ<�>��eenq���ҵ Tf�ݿ�������B1ߟ��;�ۅ�n�݃�Vt�"fm����� �]<�(E������V���y����BsކR�s��L��VM�������:׀���� �# >���[r����Ԏ���|?��&\����6���#`H�>�ۤ0�%���ș�~�İ>����v��s�©yo#�p��h฼.�?x��{W��>���|�#{/��!3ȡ� !�,:�k=�K�,	S�$�Z�5�K-7R1x5���U� ��ki��c���Ш\2�Et7cY�+(�<�NV���x���-�8�bP�}	�Ufʡ�y���q5�?˴� �*ŭ횩��~JA��n�T����cٔ�N����t�Y������,Yp�3�x�#��ݛ�����{�,v�U��;8�hۏ\t欶�h˴:��PH��e�� f��
1�#���H��U�����P�&�ʂ3��怹Rm ���m�?�~��I�ͼ�S��[x�����;N3�S���]1IUC���4\,b[�	pS�g�e^wϮ¬�$Xo� (�LOF�3;�#=��R+R��#�2cg���Y���ۂ6⽸��x�����1�J�M�U��m+6I�9�֞��d��ƿ'�284�Mk������i/<h$� �#w����!��n0z�F�hȬ��e��� �F��Fsð�<Z�'��R���㨦�:��N=��b���\��Ŝ��?	����{V$�8�U}�������|Wr�y�	X��#0��b�ᩤ|2ֹF;�Q7�R��N{Ux���\�8m��X��[�c#9��4h
���{�;z���@��2�' �5�C�����֬> �T�p�M1X�� �}�eO�{pj�hɱCyd��݌`~5�\j�M trm��C�+�1)F��M�#�	3�*H w�|~�ݷ�3��ߚ��^���W+��3�3O� ����C���<�ӹH��m���=�J������HYc��8�-�ׯ#���{��^��w�����ڱU����+�~�W��M�<�\�ڪ]h�ںe��WY��RM>�$��v�m�~9�s^K.�5�e�c�6%^�t��y%�q�GOzo�m�@��n�^{%��� ���<b�;˕��O����\Gp�I�\m_Z��\�dT��5���KOLU�O����T���&���4}J;Kp�
��V�a id�X��=+��}Ze��� Qkww�3}�R]����[L�` u�j� �l��� *��ݾvc�V���3�N(~#��'�3x��A2/l� �_qE�����k��'���!x��&�O�~���1�q�sn������,Y�O3�5n�u��o>��i�{w�&���P�"��� �Udm��Iq�iɤ��*�G��@��N|�����d�7�/����L��{�vj�0�{W�x�1�z�,�sn8�Z�]��E�±�Q�N��$f�ǵF���# ���S�TH�w��DlL�暼I�����<�=���=�:���ۺ���M���a�~��/��#�Vd�.�8�k�jBta�pN��g=��|'5h�-� �*{z�E��[Ps�YV��}�(��rq[��	mJ��:VOb�|a��&��3�U\�ך�%B��S��k��#0kq�psӽx� yc=���'%M�Ve��G�J�IhrNrJ��L��O%mӮ+S2�㷦�� kgEe�֋��̎�5\~� ���S����LyZ�έ$��`-H�?��sK�ԡ��M�`8�Zf�u-�s�͵F��zM[_��>E�e��r�S�c���j��88��Nj|y)rОF�N:�Y��Ⱦ�K�������.�w6�lW�x��rM9I�XJ)����hsHb?@X�$����&���r+����I�E��NT����'�U�6��7U���r����Vq�l�$��^M�i���(vYQ�6쯯�Υ��[]b�8����������cU�~b����ǡ�^��4��'�v�Y��
  �9o����{������;�� !�y���U`}�Q����`ubKZ��3Y�̼\���y�x�ec��@ V�Z�-�x�U\�ކ��L锑�u���\���rǦy���X[��o`>��kkǈ�� �U<�Hg��>���~5�4v� 6X*�z���U��>1��>�{����/C�����-	A'�9�)�� $u�;�j���v����8=}�f��޽iG Q�w�8;z��S��rG�C@p �1��jN�n���CG�9�ZV���?� 3![8��ӗÆϱ�hU�ǿ=)ָ��*���ǽ #FW�f�<q֣�8�V/U<̎F>�]�O\RaH`3���m���SVDe Ɔ�g<��!�Os��O���n���[��%���Q�m=u]Z���`�z�7��#��u�� 	�h��,�4����I5�(#��t���]� ���W���P�׌�I��3IlO7�$�Ȇ"@<~u�'�n5=��<�۹�Z�ltk���)�0��~2�����O���[�ۮ�r1�����K�����O	�妍p3�s"�?�ӥ{_��^�O��?݁���7m�q�OJ넝�i�����+&��o����:�cb�pP ��|rͣ���u�u�o;L#��\��Rw{�GD>�V���ᗷ����_k�gof��/OjӶ���ռ�$D@�\�NO�t�"G�x�;��DI?է�G�I7&��!���'P�-��<�UdV^�##<א��p��*��㗍a��i-�(����.2F{L��GR�����L9V+��\V����U��#R���+��O���2Mu�c��_؍cT�,�G�����i�$'�1��2���(fѴ�0��c�|>��m�Չ�1Kc��ֲM#g�&���'�l����)�ɬ5F�v#�f��M����M��0%X���;W�� ;/^Ek�Hc@F:q��}�w���R���5=�0+忎���~ЁF�s�@�)K]H��Cϴ�ۨG��b:��s� �� �W�����D�;T�qǵ}3���]xnٷ�3F��ª��;$c������� ��k�6C-����䵻e|�u�<?�Ekyz����~���W=K�O����X�x��ɏ^�W�3��x"�Y��	��(l�����5σ����
 �k����׎4� 9i<�L���2?:��̫w>C�6�I��C�?/�P��y�-A���'q?�x�PVe��	O���?:I&���ѻ��F��±�����~=E5�F�f
A;�*�1YKq���վ �n��څ�Z�*~_NyZ��Y��Rz��׸��?�߇�Nڄe��w�aY9+#j{��i�?�z��#�l�al�6玕񟍬%��u� �s�F0G>�����}�Cgq�o�Ҭ\�=��M&�5����qs$��8,rRk
Q�w:*M�6g<���#8�pYCm?Z���tc<��Ȼ�6�>�+��+�����W��S�#b�+u�y4HN܎s@	�h�#9 �5�|��I.##�ǀ+�<+l�:�)"dn����:��¾*�~�]�������̬J�Ҹ�I�K�c�t~)�wu�;+h�Xg�e!p�����UץK���98�nX�����'ͮ_������<"+pO��
��s�+y �������X��T���Ě�7��n|tǵy���*&�mB���}����m`Z�5�ܪw��9�<�R_۝��X�S���ڶ���2�H���7�r�`v�⵴�'��Kc�[�F;� *ʻ��u2�;wq���W��;��Z�v�̱��:���u��q�:��߂?�2�^��V����Z�0�BG
2x�U�ջE�Y��c��u���Z^6����._i@XXHB�̄ot�c���� �ֺO��x��ÆL�㓟s�\�7���Э� 	t�� �~���ҩx���~����ʞ!�0��8�6ie�x�Ȗ8�e�c��:ֶ�c��k0E����~�4�bv�󂩎�ً) ����M���`NP3��\���PdN_'�n�^���֕eU�s��Kz�Z�{��� �V�0�o�*��#���[1�'��'�ˤi�e�#�:�A��sZ��q����C�v>�⸋�!�YX��rO��M��Ǡ��:Ϊ-UYٯMվ�i����*l� <g�=��&�i��y�#.:�"�����A���E������6�5:���|���xwķ�|lD�D,z5WI�H5to���]G�+������k��Q��R9�t?���G�^	o�(�f�@>��oΨ��T��Ip�c8�Z��|6����p7�\j��K(�#��NʒvH�� �`#��o���+����k�D�J���I�RI¸8�<3i�xr"c�c���2Mv��z����Kma�@� �e���gQ���5�4�I�9ڧ���/�³��|��5��=�_3j�9��ڤ���oL�RjK_1��5^1���^�=�Ѱ��m;�J���*|�۞s@62��雾l{��Vp���� ���U��1��
p�*�A������=������6u����֚�w�  �JE������]��#��:&]��z���2.��^j���*�-O3�#ҫ����n��jޞ��z����sUy���GF$����x��8������ ��u��$+n����9��9�3��<��|����;�m� �U ���ϥTOJ��=GJ�ٻ��Ӽ�냜��(����⧐v�=� *��p؉d���W='P����y�+�ُ�~�}�ۭSX�*�,�� i�Re.T|�u⋗�N6c���$���23�����aa��Kԭl��xv���s�J��<󞔙I��� b��z�H���t��>�Q��zR�� ����9$�z�^����>@nP8��5�R.��|�.�	��6G��R���"u��<�q���K6�y裔 �?�^�������my�$!�����A��5/	�7�6:L�D��<�ܜڝ��������XԠo.}��>`i��}��c����Y�N�Ռ:��K��{�|Թ+�)2׼�[��&[��z�Һ��#]鱈7�p9�GNd���R��k���z��=J����$�f$��U~�t�!`;����;w���&����Hcf����c�@�J���M���%C�A	�z������>$7ct1�|A־��%�V��â�n�x�v��{�V��r����'����Y!�v0����RY@V99��k�� i�?F��`����U�g8��\F9�u$�� <T�b֤��ߟq�횄�ˀ�������Ryc�1�ӎ��-
�\>�y$�~�B�/�Eg+/f9��WU�o�i�YYI����6�0?�5���|��?N����K�g��q���Z�d�j:���7�l�U�<M�ҧ���x�$�:��
}+��Cྒ�:彲$��!T@�3���� ����M;��5�v�x�V��^*�Q����1�*��g0�z�£׸��T}���61��������G�<	&�+s4x�"�;��|�@�Z��yh�/�P:��C.2�*�t~b9�{UX�U<���$Y/0��BB����g�oj�A���_\,м�� (&�'�m��Ʋ�Qy*��������Ώ�h�ڡ�sG�;L3�����|E�E�M���hiN��[{=eS���2۩I�/�y�M��\[������ {��E�;m�3���ج�#4}0I�?_\/�_�:z3�j&��Xdv�C���`���_����=����{/	j�帞��IQ��A��f�O���_�VR�4�U���$��_b�h^�Y��F���ΑW-�#�)����S����u+�]B�HS�w!r;�W�R66��q�lt�_S�њǅd��Zt���k22;��{���|;�f��23�M��r�w�&��nG�_�^Ӵ�5�ES���m��5�Ң�9-�޿�-��ZLa6��?�lI�5c��#%���`��=jX|?�Mo�������l~`׾~�?��kڶ��kxgd
�n~����Ʊ�O�O�4��8�*Hj�q�V����Gd~k6�,sK��N
���ۥ+_<�X;�׮~�^�|'� ��Cʚ.v�c�~5�_E)S�� �Y�\��}*�r���q�Pw��v���g� j�B9YUT��־���>	�� ���F��ɉ#n@Q�z��ǘKS�+�Q��9�`�8�e�i'�֗���|X#<��g�¾��!�{M$Gpꍷk��� c�Z���জ|y��j%�m[��vܱ����5'��h^)�-���mf�`��������$�}ו4e8	�� J���/�:N�'���1 �D �z��u�>��!|n(���r�\`�� Z\��s��kw���.�C�_V�um|˫ih�!� ��~���V�G½�F��[���w�S�g�\���3X��,6�}" ʛH]���=>TO=������C=����N�^կ�o����5�^��-���'��MU�[���U��	���ל|^���W���]̾Zn^�ׁ� ��
z�xoC�|Iu�Zڼ�H
x��e/��[D�"ƣ$��_u��|�����
��'�ie�������_���dԵ[+H�n��l]�=p�z9:�����V{[��h�9#;9��󫡾`G�����������m"(���v�6�᭣4I'!�_����2�����,O�o�@x�����W,��w��S'�u1�����}�
~�;q\R���Cpŀ�Z|0��	=-¬x���PB�{���lr)w8���\~uLA�z ��U��MX�`i�>����+�a݌i��ϧ#�a�'5�?�k/]�R����2��@'9���:���id DN�zg�����r��<q�	8�p��ԭ�1�
�
�s�?LBlf�p����4w �2H�SC Y�5H�$�sd
@wci<IjI��\���o��
 ́�|]����_8U5�V�+��# zq\Ғ���|%���m�a�h�̸qc,H�yݶ����3ǯ��ı֡yl��r�]�i����v�k������}Jcq݈݇ן��W�.3����%�r[��xWL�QҦ�ܶ��R
�-�9�=?�+����"��u��NR�RG-k_B��T�s�3ڻ\�{y=���� h�ӦGO�vV��7L�+����q��T���Oee��sQ�i���uU^����:���pm|�%�o���kw�������+�kP@^�:Xׇ�?\�3.�Z��	,c�S��v�qp��w��ҨGo��S��zg�#�S�]C��44��isJ$|�bUUHǮOz��j��HO��D�����w>��������m7�WZ~���G���f��wwgU�G�0r2I�5���8#��o�(*<��H���s=�m/�VJQP�`;=��_]֛W�B�ߦ?Ʃ�\��
=׽<B9�����MF+P�z[���'�>��x:5�I�x����*�WnY�xS޻ت�O��*g�<c�T��� 4k�_*�w{Jg���ܡVHrv���MO��������K�E(����>���eHX�_�ҐX�w*���R��|Ƣ��d�G��?v����8ۚU�� ���v��H�*�?�8� ��摛nK�4����;��7��$����t�{���G�ρ�
݇����s�'Sԍ���W�_�/���y�$$ Ì��k�_�7"(���q-;+�Z����B�a�O*2b6���צi�l�C\�$�����?f7���*�z���jJ�E�F$���7�K#m�_nG9U?���A�Zg-����W�lz4~�'ދ����nqY��]��s~ȶ�����=S�/���[Ř&�@�\�}k�{I���B��!w��ۃ #�P3��wڜΰ[�	㊱u�[]�LQڒ���O��*շ�0H$r+Э��B��ҎN��g��� �>��λ����^|��k�(��-ۂ�g��}��tXǖ���p+��O&����u[}�C�H����b�d��i")bW���+�_^ҭ���D�#����Z� f�E��5���G�^�W�x}�����+��~�w�fX�sҾ�m6�&S�(�ҽW�:}���eE��
\�d��ŗ߳��yn�O-���T�����Q�eL�y!��Wݱ�����c�6��	5|�Rg�����b��W��Ƀ��cIv����(���Mu�O3@��rۗh��_����� Ҹ� i�ѱ&1��=Z����ٮ�G�	�Yn�l���^���R�#��(�6y
+��:3#�L��|7o��Ju�Iْ�����uO�ƍ��T���OZmR[�LA�w��������;F}1W�{y|��ݟ#O�5�M��^4����{W?�[�W���a+ƻ[,3�ƾ�[X���ǵA{j� c׊~�nN��e� �w{��A��`�88��F�o��p��\F�g�_dx�i�G�s�V0�9E�ڳm R@�����?x�V����x�@�X��hM����Ye!�,��Ҿ��E�y��~u֨^�A�����g���!4��3���*����n� ����\/�p�[��?�~U�2��Tgަ[h�;G�JӒ$ݟ	���p���.%��>�w��$ҬR�ݰ<��u�\f���:�P��oEv26���(�ԝ������Y,�rq�8�?Ʊ�_ًO�V�;� �o��s�q^[�Qi3�*	�N�w��禩f�:���g1�!Eb:���M�.���mb�����~ �爵"';������ƙoⴒ�c`Q�:pO�˖7����_���L�-��IA°ݟq\�</u��v�J��i��I
�6p9 ~_��_�� �f�s��m�[�<�[��ڱ5�ٗH�G�5]V�仝�e�	$���\��g���E�pF�9����[�z�}�$v���[�W�g��d��z��RY�#�(:{�v>hl�@� tV��'C�a|/��o��hߟ�<�R
j���)<�5��� 
@-���?���.�֬�`�\qK���?+<c+x��ق�<�X��< {g��zּ?%��0H��\y��FN;��q������Q��$���*����W���0ݘ���c5��Ε4�ʏ�aӢ�C�,�����W?}��uu0��W;��k��� ���k�G�ϩ5��<hRG!ke2H0�ڎNc>t~w�z	��%�Xmo�2�oj�ۦ���
�q��/��}�����6��ThX���j�~�{�4K���Z=�.�O�{�f��]�W�ei���W�|:�2��V�~}��{( W�~0��t��$�0�~_�\���<����E?�� ��V�&�g�M�E���u-�X��}��B�s���� �^��D3Y�'
�{s��4� ٲ�V�Q� �� )XWL���ĖQ�P]3>�ǔ��<�����u_�-�h|�i��?J�J��EТԭ�$QT��{qڷ�I�=��� gA�6�U �2o��$M�L񜪷����h|;�cփc3� ֯���*�d��$���r��쟥�7l`����7{��zF���,,s]٨/�"��x�]�<`W�^�Cg���lA����i?�5X)E���jʺ>Y�,o.��%c�N�u_|;wyux��A�nt�__7����忕�� #?�t��3�h�ȩ���#�V�������C�m\Cio$�Xm�y�
�����(� �.z��{���i��wS���G#�>b�� Z��O�3�r��l�ܿ0� ����E�k��¯��/�8 s�ղ��[�q\ȟ4����z�>
�4�%Ln��>�cP�eo.���|���"�]�%%&|ץ�M5�X�$g�*��t�����?#�?�}���Ι�_��gLm����]v��_F��%{X�/L �[����^'�����}�NN�y��:�4�+y�v�Q_���ѧ����WҲ��x��bc����'��m�%����������ẟ��m*�0&��T�nh��~���	С���;�v�s�7�#���2�,m��p"�\����б��y����q�Z.�.>��J�O������x�H��28�_9Xۢ�bC�f�>�h�]=� ��C�j�?
f��R@ʹ�x�V��e�gˌ�ֳ�	��x��*���p�5��=�:��.	$/p?ϽG"˷�=;����x�c�?=A���[���	�zR���g�F)3�85"(��ր^���{Te^iF��<� �<b�7���O� UX�vé,������R[�;����� �t#���q�V r���K/$��<PN���6�p�ҥ�@w�d~"�5Z9�`�yk��L��io#��P�Z�`	��8�Җi�����̡@�PN�bZQ�+��'*<��!���?��z���;}B�<�$}�a���o��G���J����PHS�� zַ���#B��LO,pHW� �z
����Z�P�o.!���2�q�88ϽtZ����>�ԧֵ�˦/=��v'��������GŐ�����+61��Z�'׭s�����~?�����!�i����֝�94���L�P�~���'�H�2TmP0q���W�~/�@��o�� Mm���z���U���?���[�L�A`��$� Z�Ms�~*���/.#���Fߜ�s��L�Dv9�ny��o5�,�@������$s�W�V��#F��`+�Oڳⵧ���G�*�#쇀����m�9����k�fտ���/�V~�q�)l�t��9��7�w��n*J%����`a�5~��X'�����ԟ�����X�V8_l�'�
��i>���Z\*��62����:W�_��Ĥ�>�a��#b{z�� ���%���!w�.�{8�R� ��5�Ni^������5+�d��m���a�|����W���_-<u������]z 3��ׄ�6��0j$�7�vW%NE#1�ǧZ\C|ˁ��e��-F��B 	F�+c���p:��>�Ι� ��1�iD\��ֿ;���o���� 2�{�����ʾ�����xv/�S�nVa�q����ls�M����t�7���Q@Dg9?.pzq�M|i�2���b�C'��C�x�>�½������G���� F�����?�ޱ���K��1�2��䟡�(��N>�����7\|F��k��Emib�:����_x�g���"o���W޿�핥��	��ހ��{s ��'%AS�F>��������څи���c�˜�8��uί}M���rn��1���5%�>L%��� g�D�P�N9>����ppF�Gh��_؟K����˨\�b[w�!����^_�D���\�����1�h��g�^�8��˟`�Η� ��!9�ʌ>��^��|�m>�Q�Kw��ZG�$�q�ֺ.r���yo�G�k�'ŚпS���q�Ia�}k��/�����y>��۸����S��і�<C�̬��H̿�嘁��+���������h���#y�����~�����������{6��у�r� ?ҽ��z��
���]֦Юŏ$�
��9����O�B�W�4� ��I��d�ϧJ�}�φ>$Cm&�$n�c����ZD�k�k��5���[���l[�L��z1�+��t����Py5���A�K�����|?,/s4~Z�8b�I8P=��+�+�Q4(�A�fN��8�����n�qu����S�{�=��%�����a����O���q#�޹gc���T:��n�վL���ǽR,���N��hzڪ<af�	`u� ?�v:/���|M���7f\�!����ο�_�;?
ܛ=K�vs�܏����_bxG�G�<?�-��"��F>�իz&cmϚ?n]=-|u����О\|��)���k��T�^28��]��>(G�W��X��;kue�\�9�����
�.I� �w4��H����;�O|��Џ��a�e	&����ۇP�q����0X%iw�7y�+��?�ݞ��	�@��km��`{��ֱv	&ѕ�j7���+�ie��̄�zS^ݮk6^�˨iP(��AI�ݽ=��������~�����b̠� ���~U�o�-?�_�ˢDp�*9�d_z�X�+�ߴ_�>�<j5[�6��>bXn<��w�|1�����L?e�`� �-���#�]^����V0Nu<���d�W�|^��-����v�a+I��_�-����t�ϣ�.M�	^h�>������]�������M:I�B���[��U��|
͵���mz;[�g��N�H�B�G�f�?�c���5�LӴ�K��GxՑxc���KA(��g��iw��:t>!��r�.�ǜ`p�O�zW�<?�|K�%���N[1"�����H ���>�a�BxN�¶�X0���p�8�Y�7�a�����7�D�peE�=Gj\�0�l�/�k� �F�iʃ�^��� �oX�׍�ŚV�<bE�X�7�l��O~�^|�!�f�XX�� d��+|^��O��.e�.0���4���sNOu����#����0# <�O'����W�B�6`�һ�^=_�_nu�ceT
G�q��ª��k>gsH��Gݟ�N�?��s���� #_}	F�s���	����L��o��Wޑ��:����%��[$���h�+3q�c|����$`�${Vd���F84��nTP���Z;B��H����"�c�1A��
y��g�z�`~6i��xޠ^küxf���#d)9��^�gp�̭����5Է�!�iz�m>��B&_[��ԃ�ލ�?)ɧI=�ML>l� El7�Sff���p:�I7�K�S�"�����`^�|O6�:<gN{תi?���٤1�(�XdW���uߏ��}: ߾m�� ����w�o�����W�4����`!��;Trٚ�;hzM�큫B�pA���+��n-CL�����D�ͽ��� �W�Qxp�H�!��ʽ��_�'ď��ܴs¹Fy�	��j;�9=���s���� hH��)m����Pm� H�8#�������'�_�,��%��+�+�n�`����Y��~i�5��� 
�ۡ;ٙ�s�Ȁd�j�4���A��{�_�Jo[�x��p@9�~2~�s�GL}CLa��b�=��M�&���0�#>8ʂi���wL��}���|)������{�; ��+����_|gg��-���T�6�՗5������b�;��M�B*�C�ѣ�v�,�1Q,�����.8�h���Է�I��2`c�Ҭ���3�~pq����z���X�n59�eTm�ws�9���ao�]@Y���(㓻���^�ޱ��N<�Ͽj]����펔��x�!��Kҥ��s �˜�p2k�#q!H�Ts�m{��A���"�����?je(�1��~� ~��[����B��a�A�\�]��>ivzm�[[~�D��)�?:���)�^�ϙc��}���~�1���.���Ļ�E���Ñ�� ֮z�R��8�$�Z�ccw���`��|������!	���ĝþz�_������V��6�Yێ�����!�k�[�x���#�0ˌ��zgҰ�F���b�|��o.��I$�9��Qx�`&�p��q��⽳����m}���QNw)@~]�ʸ�K�����}��#G�Q����K(8����2V<�6*��}�qN�La�$+� �uZ~����+R��Oj��3��y �0Y��DHI	9��r3@�!|�Č�M#~�v��\q��W$ʃn��T�xS�>�P3��Re]� i�܍��t�W�3���W��T��E��T��� ���P�?:$�*ڝ4w̷H%O����{�+���0$|µ�۷s`g��*��8oJ�[|�I#՝g6�S��l�Dw����<�Z�3M 
�\��g�6�y�z�֋����1X���E¯�i���o���5�#~3��"��{n�n+ºi��+�{z�W[;x�����{��x�;S�����U��J~__�U�SZ�[����z��D����[�o:2�W;}����0k)�5�亅�,��d���1�p�uҳ�<'����u�-����09�jQ�����ێ�դ��R�;Tʻ{�ĕ�����W)�S$�Ȯѓ<�F�f&RO�TJ7yV�jac��Uۻx�9����A3�U��}��L�:˕�gITzՔ�g��HʎzՐ����],+�QO���娮���(5��O! g<W%�Fѫ�0k�uM7{k�մ��qߊ����g��d��]�s�����p��8�<�[v�,�zw��ߍ�/5mfR�V$7��Z�c��2Z6cĄw�Ҳ�Un��7rF*�<qU�D�M-��[z	-O!�Ѻ�<�י��0-����}9�Z�<C1=y�y7�>k[ÌaY�!Q���z�{��P�� -�\7o�� ����+k4� �bB�Pp�=���kD� �E��q�:Lg���/�JK(|ap��R��K�	��W]^:r���߳E���8������$`�c��k�L��N?���h� �l�d�	�ǹ�U��EeO�C����
��*t��5V9P`f�G2�w�.��/���Kg��ȧ� '9�*Ӎ���N�c�u�%��@FFk���H�a����E��� 2��/k��t�ѝ�9��E/���&�Xt�� ׯP��[h<���L{MIة��Ϛ��mz*��L��u��v��(+���Z+�0�mr,q�,�bf{��yM֞�݊���Ė���Lg"��m�eqYKq����<�8�Lׯ�N�I�ڷ9�^}�h��#���z��,���?�ʦ2����,Gk�95*�?tъe�ޤ�~R@��c+-f�O@k��g`��gҽi�[9����.��\����&R<���fz���'�!ݮF��-�]%��섄�|'��z�3�0"��w4������� g�SGl9�in3�*�OA��^f%%��{U]b�d�p}��砪Z�%�� O���z}�L�95���a�qڽR�N�;pr{W'�im��ֹ_�n���^�˻<}���67sҸ� ���dA�=y��;��Z���3�u/�RG�NXF��ޫGp���aq���u#+h��ߚ�"[/���9C����:�~"c���H�� ֭"OS����>�� ��<�9�~U��,��79#q�W����/|��1�oo�?�|��h1�R[9�1L$Uwef\c���k������s��?
F���@�����Q�f��!��sSl<�F�X)�4 ӎ�`���?/Ε�l��FG�i�v�
@'O����Rp��A��Zk7�@�2��������T�S4�'̣��n�T1���Χ�����0&xe䀧�Jz���X*��*W�{S�Z*>U�<�:xziv������ۥ��
B��YɮK��m8��ҫ\�I{ w|�0;��C�'9��LX��G�:R*�c�<�8�2�!Դ���HA� �gbOk���G�Vj��'�+W�;�Y�6����N��FN:�h��I��#4�u�({Ѹg=?�'>��@�2�}�á�ܚ����ܨ�o��V旨�h�����I���RMK��	��jA��Ԟ*Ɵ`�ٓ�ӵ0&�`2:��
���PO2��j(#�?�]��[x|���|��f���`� J`3R�]�{
�;7%��<ǌ��B���) �p�X��sS6���ϴHS�&�f��s���Ï�/�l��y�=Fȧ~�$��$����?Ά��x?CH��Ͼh��>٤�q�r�e���6�#��ڐ
��)�#��%�ݬ�G4ʝ���g��Uc�*卑�#�*�MP�-�֩p�s#H��[88����J�Ahv��@�i����p�a<� �Vjf}�K�� ��-GI$���B����?6�<��=I�w.�����T-��s��4�/���\�����oc^KJ�K��v�gSӷJ��j1����p�:ri��MSW�·ʵ��ud�Ƕk+����My)�<��?J�53��L�Nr���_��Z���o9q�?�;���A,�9 ӑC`��2{R�g��1Ȼ��Ϙ��x�Z���J#��NP��O֡���5�����$z�/�h�9j�@��i�9#��5�E����"y��\���z�Y:f�ڔ�_\��Y�o�������w���x�վ���F�������������d��ܑ�H���0ª����8�� �$0���q��S,c
�rE����;*�A�<U����E\s���x^z�b����y�4�v�Xw}y�Ү���9�<S1���T��zu�P1Ll���nR99#ڐB6�,�q��"�\e3�_�����;�rIOO�Ib����j[o0lq+�۾�r9��|�G�S����?�1Xw�.de&BH9����s�f�;��^y9��A��w���\1a����Qv"D�f�/����?΢�'2���F�s���i�� =���&�$e�5��2�X��'�՜ewu"��6�H���H��y��
��?�O�qF���a#�|�w�� Z��݌;J�񨣋p8 �j�q�����P��>�� �wƭ���'�$��	���r.�@k��'�m� ^�)� ��Q�@����I�����vu�%�ǯz�T��T0�����}���=)XE%;''毻nU��r}j�yh�OjhpU����q�,�-�F��o�������Lŭ؂R�^��Et�Mďϭ{e�����8=9�^���;�O�NX�+h�{�n�O��6�4�����8�S�����Fc��9�K%i�~m����w 3�O��[<�翵0>���m����Č㌃\G흲��֢a9��A���~|�^M៊�υ��ͣ џ��p}zb�<A��K�Z�Ƨ3M<�]�N��8�k�j]���lv>�-:+�w"�G� c+]/L���ّ#XX��R?����K�-�UF{�_���*������(e]�ќq��#·��q�X^X�|K�?��<��;Y:6]�.��0�οwP�� .�0ǥs���w�^I4�����=O^�M�uC�*�ߚ��X�O[���~/h����"��@�����Q|`�t����̒^�,AOs�&�>��j�h�y?�z�P�5e���2J�c�4Is rw��s���[=3�f��@$���]��.��q�{�
�k먼Q�J�hΓF@���_�6'@���pO�}��=b�h���B {�KttB�?������.V�fp�0rs^m8��\��NU�g����;=?E��0�$C;>�?Q���Z�*�l�3��A�g=Ϧ��\��t[�>�L���*�ֽ5��oi�$@��X)�5�W��;���?��ڿ	��J0�����Gm���h|�����#st���pȧ���=��^�dw�1#9�?J� ��-���4V��2+9�>�
�q���S�R}��q�7�kZN�΢��G���~
�]��@Y����5�_��#2�hd�$� �ȯ�<�P.r���?�~�g�����,��x5�[G[ғ~��� <#���m���v�ݏ�_?\� ��:�<�v���+�]Mo�|%����"��� ����_��B��®޸oQ���N��ȩV{��	������1{���
���s?�!y��ȇ=�_�^$�J������� ����:tQ<J��Nx����:���d~��|Q-�ݫ��p0=���� ��<Uo�O��Z��b)!��z����}}��2��S�=�A������d. �s_|@��?]~����l#��?:T��
�害BAG�B�����Z���I>��J��\y�
#��]9]v�gf���  ���V`w�4�2�����?�k(N�!5�xW�rx�Y����{M��b����$�ڽO�s�������eR��(;�@XP\O�?g��ǁld�u?�A��� 
�=?G��f$1������Q�yQ�;�ڷ����VRN�s���>72V���6��J�c�V�
0=���+CC���ۼ-�}x��f�9���Ia#��e5rU\�Т;�6�np�U�\�1[�
�@�8�5�9�S&�LVb?qSyG��\h��S1��C+�㎴�z�Ҟ�w<Ҳ��₈�0��U�۸���}9�e�>��$S�W$Q��m��#�֞zgo=1E�4.ե�~4�����.��=Gj`4�I�Ts(���*��#�)�EF�_J�m�2@��F�i�G�
�t��>��3��Mc�<�$]����Z3��J��� �T2|�y�4B���5�jX30���Be��N��_\m�U�W<��}�.��o7m�5��*�9"�4�� q:b�!��#�ҩGBY���db�ŧ�nFktB9���, �Dc������?�;淄��Wg4;q�k��|h�#$�Xh���B�ˀ}>��8`����FQ��Q�ϔ���^Q�ق�\��w#��T�p>��ǉ5B1�1�9�I���Hx�V{�0��9\� �q��T�F��|�}{נ|
�<�4�挴^j䞜��s����5�\�k�g�u];�I-癲Vg�ݸ��_[4�������7g�$k��V�2:�%��p
���9��>���y	�V�.2kW�KC��`T-���� �4ԛv+�Z�g����ZԵq&EQ��$q��cl�oj�(ɏ��s����Ḙ0��շ_�5���犷M�^�E[)���ҵ�jp~�pہ�4�0;`P��cM��Ӷ��s���rs�җ`eȦuշ��0�[�X��:n�Mn1I�8�<3��q޶����"Q����q� ~�IPGA�M$��F20 �v�J�g��=��:��ZH�E?/Ҳ��6쌊�e�^}y���<� r��j���,�>��"A�o,gS|�����}
�o�d�̅x��O�Ȥ�$���Ҡ�@�GN1V�\1���"�����X���k��lX�y���Q\F�5���9���YI#H��ɍ�8sWcfU�K��l[�ٷ���i�
�̨e=y��fS����]%{�=��=8�*�X��g1�z����F�r��d����4��|B�6�*�?.�[A4C���Ĩ���l2��В<�u�~f�:na�nM}q�R1�u�1��@_%i�X�s�F;�uȭL��+���B�s��sP�e c��W/T-�'�j���ノ�L��`��p=�P6�d�q�/rx��p?u����<�&��yy�?�n�I�����)�H���9��R���F �;R��Y��Mۻ>�?�^�Մ�'���郚@x�>��1����`q�( ��o��K�h����RF;
2{qB��&M .M!����ځ���o9<Q�.A8�h�)���}�A�{P!~a�ri���֤����{)� �{T[Dm�� ��Lb����_���1㸤������ml�f��5C.�Q�z5��q�je�Ǔ�?���6���$���i�������C}t�v�z
K��;
8P*`i� 7pA�mbyp����c����5j�ՐI��[��DA_j F��N��M��n� ��}*�32�{��f;�$��=(x�ƽ���U��A_��g�_�y����|r�4�-�_���D(
� �
�Vc��n �e���4�jyI�~�ҥ��c�� 2z�c�Vj�v�͖���1����� <�#��o��I�����$� x��2�P3��i�ȋ�2ZA'���W4��`�mN:��t�r����&��Z�����T�8�� 8�A�jig�,n�=�	|ٜ4���R��'�!$�v��[N���L��+�����x�^��$�~lt�Yv��
���jmUڣ���MҥԮ� ��sϡ��j�������N0ϰ�h���E��So�61�kO�%ԤwN�[�8� 4m��������n�����RkZ��a�y��(=kVL`��X�+.�c��֔Z� �~��n0�0=��Tk�|� q�Ƨ�֚���*�x��S�m��9��$xd�$:T�1����8����4�To�q�S���=}�H��t�Rc��VP:�\�[�~\���֧*rۺチK7�PcҤqr8�@���vpq�֜���piT�B23�����a�'nѐ3�3�HT�|g r1�z#R��?���)ȣjg^�{Sd�_/��E\Ǯ=������d�8�R�!G�{z�D���&��[c:pF:S��\��P=@'@)>�G�N�:3�q��,6&+��;��0H'�P*�d���N�A���M�8�H���	�����?����W�0ɋDC��+��'t�� >��T�:��l��QeW���Ξ�˞Aڦ����#=i-�̀8���U�<
���Ċ�eO S6��h��j�	r2{RC%�\.H�S�S�gJ��^g� s�W��l��"��Ľg�A��X'���u(`q�n��������Gʹ��W��n�#����[GaOr��W
{g?ʡ�,ԓ6��'ޣ�� :�0�Px�4�bܜ�ԛ~P3�ޚ��0�h�S���p��N��� :1�q�� ʬ�t�h��8��?n0	�����d�@���`s�z`��H����$C�c�;�m�+N�o�*��e��ů�BNCq�W�W��~"j�vײ�q�fnp�rG������5�֍� .r:�2���#h~	�#���4Lf$`���
Pi�FR�<����*4-n���F���t���O����~fjү���Gɻ�{1_��Rߊ�$�	���%��C�Dr$
��>����7�3 �9�� ?ҹ�����W;?��G� (,Nk��w���ĭ^��p`�b>|�}�O����Ɩ��3�� ��o��B�V�lגƪ0��1��?3[ƚ�Ԙ�ō��?g�v�G���Vz}��G#��T��׎}���S[���R[DX��wE�L�_����V�e=Ǉ�����L���rpI�_�E�J�vL��>���X�M6T��:����Tgn@^FZ���_�j�<�l���FuM�x'�_|<����y�|د��ٛ�W��+�]��yc�i$�����_��w���M�=
Y|�.Ey�� ��A_�_����*x��G�(�mo��/,��d������y��ú���.4��ZKx��"0�U�nLz�W⿊���<Y�]��&�����qYS��*rm+�>�?i9�񏛧_�}I�'EmP��@~fZ���F�.�|�s����>��x/^��WsV��љFN/C�;��5�m5����G�5��@ �����7�9_��!F����D�:�Q���U�k��C��m}����R8�䷒.d$z�_����3|{��Dj�a�������ci�ۛ�7g���M)e��hf���R��0�3�0)���ٌnϨ��-�G9�p�i��'�>��]��� �LB�[��u��_�~��X�|�<�8�x�#�W�ɹ���FpH9���K��� �}���G�"�~�Y.���Č��� ��kŷ0N�c�V�U�#�52/X���֮Ɓs�j@V8��Wa�s�ֲ&��;y��|��J��5#Ǟz`�1��Ǧڭ'V㑚��1P�{ず	 ����d�Lf���6�9��AHfӻ��ڒA�>�����T�&�3�RP�' c>��M�����r:w�F�����Noʣ�,J]ކ����I�u���sJ�747�Ә�Γp
)��=�#S��E��N�0:Ԁ�Le�AbrOJf�^��7��U��Ն`GZ��y�S#T`!p:�?��~lνXa�g��6ݫ�� k5�=�bz��
��2�q���
�5�j�U@�d���ж3e���3NٓI�z����ALV*����'�J|�>��L~R:W����qȤƷ<��w'nOZ��7�T7�#�W�����k�~$H#�s�Y��5�G��[r�����C]W����V�!�ν;u�<W��<I�6�4��~��j����m}�߼��2A����j��~��e����>��sļ��?�X��i���o�^���½)�gl*�"� >k���ہ�\���^�u�������r��wM�a�U �8�k����x̀���*�w�9-�nJ�o�rj���8��]�tm�<�V���k��$с�֬B������A�U��}j�X���D�
+���n���5+��)�A
 ��Ӝ�(l�9���ޛ���ܯ��� ��Ga�'N��֙�R*{/Ozc.��4 �1�?���Zs�^�ɦ� �b��~4֏�=i�z�nۑ֝�a�F�_z����lz�� #bqU�ld㊱���P�<qLZ���b��6�n[��W�k-�3��^g����ް����xv3%�q���]B�q�t�/��=z����q����X���%9�*�dR:�&�e�B�W�|B]�2���^�p�y���ۧL��i7����� �wQ\�*��?�ƾE�� 8]���f������7�18/� ���|�g�<���q�?�Z �}�ϵW�P1��U��7\�y�FH
�x���b��͜�>���['�~o�&�e�*�'qB0@�@��1-�#�;pG��������>_M�Cc'c#���y4�����֝�T��������ǵ!�h���B��jy���$z�֪��}ޔ��<w4I�Jf6��h�$S�=8�9�1�?_J\�9��?���ņ�M$m
	"�O'�hw�����1�G����
����F��w�Y>Q��o��k��Ko�FI��:V^ܻ��ݷ��ѣ*ex��-�e��P�0���� S���u����^�c���k�����j�$�)�JV��dg���C���:��
�m��Ş�yt�I�w�;TS�4�cmD���c �}itq%*��Z�FK8X�n�Ҡ;-W��Q�I3��x����6Cg׵G��F}��Ozw,I�b��8�9��)��ӯJQ��� RwCJXn��-��~([wf'�h�7�K#m�44L2q�H�[���h&�Ƭ͸|��j��n:���3���*�,B��j��3�~�wN�Z�`�mA�Z�g��[�s�Y����?*7�IPԖ�|�M��8$������̒��-��'ڝffg��I����*DU�L�8$P������c8=	��y���Yw�� ~Q�c��pP��0s����*TQ��}ia�In S�</� t�]���%d_�F^���V����4ח���7��z�V<]�˂퐯Ldc�O��L��G��� ��G\w� 7�Z༑-�N ������ ?Zˎ6F�rí�c��=8����{����R��2�ho��Iׁ׶h��n��N�F�� ֦*a2H��S��<�T\8�N,W�����R��O֧R�$V(����a�叿C�T�Ϙ�޵&�<��y��з�a����M?��{U(�+���q�\g�Ӽ�V��;ҷm��N8�S�R��NJ�튉fV�\����=���v�2U�޸?�I��2G�S
F}r;�S����AS�΁؛s�#<R���)�9�������d�;i���h$zi0ǯJjǷ8w�Ş�i[�R���JUN�y��z�;�ۋ�h@���B�F\7�ՖV8�9��(eGt}�� �q�u �n�t����󯸭c/f�=*�g�	�Kx7U�r�x� ���
���1���~������-����x�M���ƣ�̀pjf,çך`U�����\c�RX��	�7J l��`R4�T�i�y�MG?����G���j�7TO?O��|�3;��>���u˥�0l�_9��.��������6�-���`�.$=7��j�M{�iI�=*����<�3�Ď3L�GZ{�I3����'��j@8��1�Le 6s�Z7p{�H `I)�>l�l��?�S�ra^�*)dy�{ b����}�q�3� �;z�������E�6��ɧ[1�m���ީ�8=�)��d���Pŏ�/4�����EkE�{�PȆ;�be9����n�h��2˕��L�U���(��P�Z��O���3�c�u	�U2B�d�Os�L�ö����_����K0~�ϵs����֥[�$�h���j-��&�%��q���D�x �Z�� 5�[��+��vyg���d��֙�eI=�|��K�/�>#�5���d����7_ֹ�[q���EH��Fi?�����l�b�T����h���F���7 ������5�ϮM~|��V��tz��� j�-b��ܱ�,%�0�}?Z壷0͖'�zU�_$�z��W�\��9����_�&��4�&�?� }v��-���\#/�]ʿ��j��+�1�=�w�y-�E���~מ-���Y��}ӾVf���ֵۿk7z���WL�9�9 �J�&��'��1@�s�8��n��Äm��8�=h�ZO���.��G|��7L�D�[j��7;��Қ?�7�>��p:�:RϷi�o�{���_�m8����߶�S�W��`.zW���l��M �N1�I'�
h���Z܍�d\~U�Y����;s�8�/�k��m��=�e�ѩ6��皻�S����1�1W�'h���Y��h�4�?/�Q�[�>X��4&\Ry�뚮��ԫ���W?$ZlVi���Ue��6��m����/��1P�i?h^�����5�%��L7E��>�<�6ŎX��	������O���(�i��S~�9��nw T�ڇ8�h�_�K��E/���:v��F�-ןLR}��� hzt���7<���>�;�I�.�-�G��/�sG0�m5�=��p:V?ڎ:��`��s��o_jA0n3Y&���t7;��(�(�� ?@����t��u�2��*�9�l~�N+ϭv��a��5����y����g�� ���=���v�Мg�� �Jя��՛n��R}9���j��cԳ֦���j�<p{S���i�I2��������=��Fk�+�p>8]ДO`�y}�\��y��h��Sֽ�PR��ڼ;⌛�������]F|?��?��<m����Ѥc}���s�r���bB<Exq����V��\)�6�W�?�]=���?�Y��O�TcӮ+�헭y/�ǟ�T�D��;C/�9�Ez�'�'����X�jʠ��Sǎ��R`V�*5�+0 �U��qJ�V � ���u�J۽������Tw�Ve��@��⋉jy��.��$�((����,�?+d��S�@' �F)�eF�Ԯ���~�6���I99�T��w�T_l]�g΋����w4�`�ި5گߵm��.���'��Q��ǃT�׻�5�@�4\v/4�����Pkͽ�����4\,h��.7u�k8^ s�>յ���;�cA�cӭ3w\�*�^s�ڕf�h��e��5���U;�y�D�y�t�I��_*0�޼�U� ���zv��g�S^e�����5�M��z_��d��u�?���������ͤǑ�x����^kx�`�&��3N�zU�NzR����9�+�>*0]6v<�^�p9=��>.�&�t�O�$�'�V��EoY�
�ҾG���&NO�đ���~#�	��nV�c؃�j��B��H�pI�8�jџB��26Fy�B�9��Y�fY��	�01�;
���y���ր#�|���������1&�rI�)��9�}�9��,���M&qLEl�q׷Z+�8�Ll1��A��Oٸ��}i���`�_ ���t�*zdc�j���Aێ��1�o���ʞy�������9��1�x��1�ıJrǻ�8�S�(f�&��*1�F70'�o�z�wnꧮz�1����9Sw'����g$���y8�zb�#�1��b��E������/��ǈ����ѷV���� �)��WĿ\����G,m��M�P�q� �V���� U�wI����V7�
���rI玿J�r��D�cӨb����J�o6����R�h���H�����9����P~Q�:Qq>���}EP�fqy����l�/\gڗ�F��O�v>�O�k֢fFUe��[Q����*�{0��r�Q-ðݵ���t��!e �3�_f|#��<;�xn���4�啷#��マJ����}WᎽq��?�+�/^#����a�U��nivq�4�I�A��ڬ��X�c�X�,j���ߝ1dq�O�UZGf8�LT�Ȱ䑖������H'�zR3$hp�9��/�u̉g�\��
������)R?�K��
�����"�n����:��'���������F�k{��'9S�SN��ŏ9G9���1�'s��qYG?�Mn۟�ߜU\�m�6ҩ�Q��I��X���`��۽8|�6��$z!� ���b1�=�/�'�杕����Hm�q���Yn3�=)��r�H�Z�6��M��F8�ʦ�f	�7ޛ&[��R������t�2� ��$6ɖݑ��?S��Ax�t�ʃ�u�*S�G~��� 
��?�YW�2�yY�T������i��� {�R��@*�j��x��{S�s�ѻҜ��G� H��Ƿ�I$�T�ǥA��df�؀;�t�ǫr})A��[�4�c�
 ��g�H����=:R,m)�jx���ls�]U���|����<��54v��y5dX��ph���q�/?N���ɂ:���;�G���׌�Q����>����d}�?/<�[ɻv�1�<�+�\rq���q��qԞsH�چ��X�߿ҝ�c9�b�F͌��#��*Ұe,H�p@�b��09�S�M�9皉���8�"�RBs��4 �c�$g$w�G�����ON5LF�zg� M�����*ڷ�y����dH��[-���~'��*y'<P5�>�� �u����tq�����>Y�+��'[��֤3� /Lq�f� �W�a�quǭp�ͺ��<�FG�֮@w.O�T��5"9^��M'̀>�_!�/A�i��+
 ����=*��qW�/�g�Q��h�ƯB`��d�����r���2�?/��+�O@#�nq��a��m��5��%I�+Jo@�����'�>�+62dmǖ�z�;
VnN<
��[���b@��]y�9�\��&�� c���"�*�h�`b�ʬ�x��s�Hk09z��K���U�r1@����K���9�Z�eY$®��}&[�E�K1��@̼n ��_%��9�����?u]vH̱yq��z�� g�&�(ecq���]t5�o��"��ѳ�����[�_2Kf�M}� ���4�q���RCw��x^h��,@����?h��[C��I����|��\�=�5�G�>��$�m�W����|5�Gvhyy��著+9&P�@�GB:u�1�x����]�1�$�� ��M�#�
��>�gi��4������L��'�� ����K���K�`c�i6��h[89�J��7|ބS?ձ ���m�'�� 1�I9�O�/қ����Niwg��:d�?�;p����{�����Oj n��x�n��>إ$m\��4(=W� 5�<t½��]m��õ��8�,H��~� �k�?f6��N��U������	��M]���m'�[�2��}+���>LJz 3��]����}�%�ѥm����5z����T���Z� � J�e�<`T��S�Q����Ԍ�)�E4M�Q�� �:�;��@�����J�~f>�CG=�?�=��ٴ�Y��ά�!���[ m����١�t�a�&��5��[��w��N�9���W9�`ۆ��oՆo��v��P͂2(�1�4��F*C�;1!s�Э��q��҅�>�r���K��JO�w<��DZE^��G(��t��⁣���C���_A�|�ytW�֓�ُ>���^�`^�;ӱ79���jH���n�ڑ����=L�{3sޝ4|W6�3ޙt��qV#��#�;�֣�x?��Fח�<ל�� �z0xˎ_��空5��6�Lq��V�9�t��Gʣ�U������+���-Õ��jP=8��=y�T�� +��	�l*λ�������I���z��R:���n���~�|����8�_>|M�y��ea�k?�2_�E`N�Im���ގOLs����� �Qy�ǘx�ޮ����
� ,p߃WO�#�\�h�����H�2���� ҽ��7�^?�-�� �Yd�o���ױC����b�qVR���C�j�l�	����Ü�*�8��
 ���j+�QRƿ�T?2��z ��f�+y���SVm����V��n"��E1��1�-��l.����/�h�R�Y����o}��n}�A�I��q��G+��sLi�kxX/Bi��#�������)�H��kut�Q�ɦ5��G+�����9&���j?��� Q���/��'�4��>ƶƚ?/=/�b�� �������T��{���ʎ�t����D.U�b�.*�C��qڤ��+d
[�+�l�9�n<F݀�ֵ������5�z��^S�Y������ڹ���� ��6<�?
�c�ڰ<:�-6NN��t����ܰ0)O�=�>�?��D��2�W��^Vm>a�<��k�n�}+�>.0\����@>T���|'}#��l�=?ϭ|{j<�&'ߏ�pk�� ���B�1���f�>�S���,� >1�*��B	>i�1P�@P��8ϥOp�d���Wc��C��R�A�=)�;���ZM�wN3��'B ���z�PF8���\��!�>�7�����2@�A���^����N�5xN��֐��� ���L�6i@=3K#|����S���?ҍ�^�c�@`:�j�����W�bc�����1�x���i���l�'֛�A9�XK6?NkB�O�c��ۚ�b�͖�þj?7{��k�	��$d9 d�� �dh��ֵ�}>�&�Y�h�h�楔�2��&q�9�ΰ̎F�~�]��߳'�,�b�[w�0���gҠ���u{�S��8��ƞ�4/���|*��Y���~��g��_Ik����.I'�}�ҡ� �Y�$��^�$c��u~�t��u�YeQ���ߐiJJ�F/�&��oX��+�bDp@iQ�؊����,�)^����XlM���������·�VF��=�Z]C�gï�j��~x1����D���?>�s���Ƞu?���Lyny����Z�u��6f�$9#�m����]�o�I?�;������{�(�9q ��v?�t��;}K\�i�pzU�K���O���{w�x��<+y��p����4}Iw��Q��m�x�ϯ5�ۋ��� �+Ʈ<_}$�Y����4����rN=E��=���u�����6��ֽS��/�������u���=\��8"�5o^2�wm�<Se��ZKnUn��	�k�B1���
H�֛������^��἞6��2#{du�\��]�6�t?��-G����X��m8�k�n�u�AVL���ʾ�ҿd�ԯ$�f8�J|�J��~�ph�^�&/�3P�_b�5=���)�'�� ��"�Z�<�,�0ʠ�8� =+��񥇈�_0�q3��W�x�+���FӰ��q�q]?_��L��s�r:\���#���V�N�з���ּ�㖗jn-�(CJ	e��:����8r�=�{π�Y·N����#tD���2](P����0U'����_X�~ʶ&2��>��+�~/x<�$q	�#�S[�#���ڹ��zr�rpC`toL�[�՝�Uɬ���t ~U�ɱ���v��Jk�"�Y�0z�d0���t4�?��FU���M2	&��Ti��QQ2d���WM�+��(�������f��n�{��T�T�*�j���z����1O��-�aGn����+���?�Ӈ��^����Ҧ�n��v���.0t��9�Chf��+�w��R�⣍��/&�Q���W9��y7�a�{S�m���?��=��\Ϩbh�~D<s�����Ac9�ds�֒V�	�:�#ե�8M��4MnV0�sSp�Mv��O���p���&I #��5��5P��;B��1�~�;�4��`��7n'hUc��+�4ٿ�Rh�k:t�M���p�`J��>_ƾ���d�/�z���;�q���� e�Ld;�}���N��g�#֯��9���X�8z�r����k�yiH�X}kr��s��2Kq׵{<0���0O���J�6Õ����?��Ձ����W�&��d`r=�}&����ҤiU�T�m��}ʲ>�<�蓺��篥`���C�$c�}ͫxvj7R��r#����,|{k�T��d�W�����!X�T]�?tt�N�a��<�Qc-��A]�wz�c�`J�Z�A��H�pNNq�S��̝6�93F��=7c�?`b�W��{
 V�ħ##��PY���pw��;{f�6���E����yȠ��_��k{{Te�H�O��vK��Y�#p�j��h�j[�$2���c��^+Y�#��ӎ�c�JAϵ���2��Հ�����y<*���J��F:���	ҁt�ne�_��} �� Z��\4c<q�q�so�A�$�槙�n'���ű�^��ͷsc��1ѻH���j�~b:T��Rs��	.rܖ��1T77�N3�*y�Sm�̕��?$�qk�C�,q�9��|�r�N[��}��Bԯ�o�1�3��_,e�eP?��w���*nX��Bs�4Ռgp��i�y�3��
�d�f�2�I����������rT26�Oq��Y�[��?h-�cV��ǚ�n�Ld�N�5̣jg<
�O���yb�z��T~��j�;C���I�5����^�)j\.и�qU�w�tӅ��3E�U%[��H��z}�� e�9��4����A�C��W��x��p=�����k�ꊻ�p>����a�p+6�WX��f�/��-���01[+��"�&��3�n+�5i������z��j�y���>���H~nv�ӥg�	�yOod_��?��yɷ�Պ>r8��k�s'M� �J�_�:�ww��m�ܟ_��FV�ɤr�t�1e2C�p>� #>�ա����A��
[�8�z>�`��`!✭��iF8�������?�q�t��~S�c� ~?JT��
p��I��H�ޑd+&Aǥ jG���i�8����{db��kM�I
9�� �K2��
����zP����{T c��c�����wX��G�@*�w֑r��ϵ=z�{zQ�F�ސ`��@$ׯ����aX��9�אc�}�0;׮��������%\q�Aq?Z���� '�Ȯ���V��c�c?"��ߴS�����ѩ�8,3۵^��\g���qW���P2u��ja��60=�\n�;�������u���l�8�7���`�ST�L}\�X��w�=8��H�Pq� ֥�[l�O�cԳE~��S��j��_Jw���Y"n8�֗h\u�K���c4���恉��c�����$ѹ��r((x"� Ȧg����I������E�8�<�:���ڐ�9�a���}i�z���&�V?�W\�"�V*E
��rMAs���X�A���q'ˊ�Nc^a`Fx5�c�*{n��y��{מ[ɏBA��k
�Tk�ar��.xz6�5��.sש�Z�5�C���?�J�@�ѷC�{����H1��v瑚�b��c�I�M�`�����>)����0k�mms/z���Z����[ �
̣�pn�E�#*]��� Z�i;��q��v�Y�:�'�w�x��d}Nj֚�6#;\c�`���[X���o��������uֽ��ӊ��;��OnI�[w=������u�P�����8��#�W��<}���hڞ��piҟ�ǽ [��v*��ԓV#]�{��&�U�9�i�F�8��nܧ֭�	��ިhcd��j:���
�Ի70�T�r�VH� (b�+��ZsdTL޹�)�1��q��p�1֔0�1ǽ 3fs���<T���8ⓨ� ����e��R7͊e 
��4���)W+ވ��ϵ 7��ڤU�Ȧ�K��<P/8��_��X({t�ׇ�g��+����.���{�U��n+�uO��@<�5�SsX���J�?�>�V�_68���]� ��cӓ���ہ[Gc'ԛ;zT�qMA����� *�H.W�g�W�|^�,�q�kצ�u��k��.�4� �N�:�[��&?�[q��l���Ɩ�픞N0s�����S�Ta�zͺ&N�k��<m���{ۜ�TGB�����ED�w��ԳaKNwt�D��鎵BF�c�޴�v���㜂p{P~QԒ)�a��FI��;�9���2�
 �����s�(p�YW��K����O�'Py'�����P���w�Si�
�k&��ry�῕H�����L��u�h8�wg����6J��4ś;�����(涴�;�Be��&�N�����X����%�קz�'�e����λw��[�9���R�9[?�>5�*Lm�A�m����|#�|;�ص]F�G�
�p	8�+�;I�����*g�-!�EEU�= ��[��Z���|Y��K�{{H���n'���X��݃f���FR<�l
�o�CV� R
rrҝǩ��8����Gl���G����>S.�=K��U� �R��5F�~�z�� �T�J⽙�׈?fcg��8o���UV����-	u�l�+�mV�-ؒ��pq�Y� p3�R������U�Uwv�]/�)[��)��+���+{�~]�Y��jw`�� ���m|�"���� �L��+k�[{s��ֽZ��n.�*�q�޶ ��@�v���d|ɫ~�6��>�v���s��4��I�ӥ}�z���E�t��?��:�g]���<����� e�S}�#ۊ�տg+H�����Rh���P�S�����4Ӱ�<����/�y[��ҽFh ��PpzW)f�ks!S��󥸐�Fy��\�Z�-c-
���u��1-�U�ہ��I-�ƶY&��/L�B)�)��Q��k��qڧ]<�L�Ux��A��T2�������5��ƭ1��VW��f[��oyr�:�JⱥͶqגq�k�_��	.<k�	`[=;�oֽ��'�M��<�=��VV�Fq�������������Y�_w����x�3M42�s��/j�	�����mm#�]Ԁrx�W�_�3��_�^�L�+��sߏJ��2�������}*H��s�ơ�F� zՋ��7����o�6Y��ڬ[�cf�I�1隅�:�t��!��%���v>Pz�M�I�*[L,Ŋ�<��L�j�H �� �Uk�WOQ�W<A�laJ������ Z�0ň�|
1�Smcڒ� qڬ&}=��љ##�'׵^��6��Ŀ1�?�oʘp��� �1S�f*H��V�hZ��Y.�Nw.H�<՛����ߊ����*��V�=�f�aX���n��^��9�N�S�:��n%ӬK◢���
�fdV7 ��fm��[�#1W'����8�O�<[�Z����>�@���ӿ�y����[,O^*o'��)e��ޣ�?�sϭr^��ȓv c<��<Ԋ�S��q�4܌g��>��I��$3Ny
��J�Ϸ���T�K!����[v;��4��4�TR��q���.' �b���~p;s�(|������M�?��$'1�
�
�{◆bռ5uq��xcg�u�,��ص>77N����WNZّ$Ih��y-�V�8�285JY03�$~Up�.3��޺	%U����(
��9�F���y8���1�������7`�Ӛ�7H����*�Q�� ��'�Z�s��,2�Rʎ�۟�OY|�\���>���f1Nx��� ���B���E������Hh�InoԹfV��SxϚ����c��V�Bςqڀ,@�W=i�!9=�=Č¦e+b1@�8O֬[&�A�w��A�T�]��g���kT��7���x�5�ū~���r{�3���'ŝ=W�:��6��p���� ��eKO�4�ܙ�]�Ei:qL������K��:ѷp'[$�v��1�
��)�ぜ�/�sJ���HUm��{�]��i�8�"�b��S�mZ�<#����N�g��C�n}5��4�|>Ӻ�����Z�3o|�O�� �~^�ix�*/�V:��Nۧ�y��ο4��r��"���g��PM�(����}k����9���u���u�]\��ctv��� b�� .:�'��qpv�S<sX�]�3��`M@�6Kg ��ؒ��{�2G\�Lef1�銋�f�;�|# e��i\�3����n�j��M�;2vn란� �iF���0���Eu	�	Q��3ހ���wGw,m��F?���L�����_�N�~�5_<��µG8�� �:�9�o��M��g��9��6��sL�J^W�^���o��=sCc��X����G��N��#)�#i���'��J�qm��sHR?��m����UD�aN[��������G>���� �<*`Y��eP3�횂����%�1R5ӫi�dq�Z�ᛕP�:sH�͖^ps� q��K7p9�\P��(�S��օ�=Im�;v�!��pzP;���l��8�[��<�m�&�1���+�� a�'�׭�̀��;$���u��Ah�p�lg$�('ר���Z������;W9�g��r~��� ?Z��Զ9楍li�0����W��T�=*�y�v�z�Q�Tun68�b���j!��T�F��MQ%���G��w�[�	皻!��Un6�R0h{��G��5J�=�8&��݀Zύ�H�gn���<R�5����7��3B�݁�5�$�Tr]"�P*����8�l�i��� �P5��?;�,3�Sd�-(���4���˜c&���S}
���=iV�-�y:v�0��� *����ҡ�Њ>��`-��_vqT�P�l� _�'���c>`'ڐ��&ե��?7��Ŭ��H��iU�H���֝�s_��3T.&�O5����eP>�B�\�?(�s���Fv�p����ُ��g9���ߊ�J�HYVU�ּ���n�V�ְ��=}n��Y�P�>�\��,�w�G��{V�A�Ov�B
�x5��B9OQ��Y�bEh��OJ�	��O"C�Q�s��;5��sN2���g'
�|a���v�ۚ��b�wֆ#�u�k1'����85�V����u��|���q����]{#ėݿ{�_��u�2($v�:��?��׬8fc���U�M�I�mV��+u�h�g��m�~�s��U��~����w|��~�g�P;~���G��{����j�Ѷ��^j�k���,�1R��=?Jc&\��s��\ԊF���w�A?8_j��Ap<�$��!�z�ӓ˙�<���q�Y��f��E�$������ y�c������2@�"��i;SJ�)�v�9�ԇ���z����@;p:�gs��Aa����a�0q�������}:�k|��8�@�<I֝��0jo��jr�s�,,���U�}������Fi<U$&�-r@���W��'�&O#5���d��Q��&[��*空5���Q�n{�ʶ��(5���m:3����@� 5�V�or���#`�J�6�O,*�A0��'��.\��ҽR^��y?�f-f䌩9��Z >k���?�$ TD��q����1� ��
@s������b�</z��17�����v�7����;�.�%c�Nq�����d~5,�|�B>e8?^�֑b�q��H�m��t�N�N2*ޣ���6ˎMG�xe��iZi$Q����)��|n�z})���8�~��j�@�K�LsUY\0���d`S���z�u�y�\�8�����5*�|�z|�?�(�vf��W��~8�aiN��噛n�������R7���.N�tX{ŏ��L��M��js�9�u�3*~#�P���� ܚ���tX���o(%	=Ny�+��z��(Pv�>�����~*�2�O��}[gp�~�h�9Fq�<��<۽��h���-lP���8J���#��Úǎig���Tq�Ri��t�GZɚZƵ��[���zWOc��od��a�r�pU�N2h���	�����^&d��V���5��_�kB���'������,Y�-��<}(���ϴ�f���zlL����i_K7�j���I&rG�h�XϾ�aU�rj�j�X�;zV����nH��r�C�dw��v+]�
O����y���U��RMM��~����HV,F���꼆0ĨҞ��-�8�Z��2@)��$b�JHld�P��8����J���a���#?�Ҩ�SE���ݑ���6l=kS��n9�cZ�y�/j�+�s����VE�]�V��ojw��Ґ�BÎ��Y�D����w=�֩����G00��:�����|<��W<`b�E�`i1��~���:�(_���LWz�Fc߹y�a+ܤp�2��1��(PT�V��Z�A���Q����:�#]9�a��s^+�\yͷ���mQ/s�?g����/J���O3�Nzי~��	���K�hԘb��g��]�S$�ܜ�~��Q2���=H�ٳ��\L�?8�o��pUN�{���)���Է��=BB�`brW�5��\ƙڬq��S]kT`�#;6?�=�1�;��X��b7j��q�c�����i6�!r�1���!*��� S�C4�s�E�
��鷞A���U�[y��YL{b�w�L��a����q�3�l���j�NO������e�FV�c��U��S���Oat�W?4tY�ƈ��H#i��U���t�֬\�+��CA���(��i�c�P2V� U���;3ģ�w��*���[ۯZd�=y�h�7F9�-��c2��y�MpA#��������ց�6��6��<㌜W�| ������
�]� �x���ھ���d�>�.�e�1'��gR�.'�^M�B9��R��ŕ�L�U����pO�V��H�j�Y�I�ӑM�fX�( /N�Y.���s�f�<�� �B�o_J	��{�dg�5NIs9 t�_���{��P��if'����=��VX���Xa1�
pj��g�8z��rOj߱��wl�@�-�i�T�������08������P�*I�f�3��Ǒ����}�Gkt��)��9'��W�ŋ����'Vʛ��ג+%/�+��8�>��Up�ȭ�]�=?���$\(!��s]���S!��]�94r�n�?Z�@�~_�G�U�����}O���P+���9��6��{⣅J�N�}b;�A���Gj�����B4=y3�n��$~�ʾ��ԛUcҾ� �y��7^N������Z�� ٪���G�s��T&?>L�&���G~��'�F�G��F8�Q�H��txn:P#c#)�o�I�C������G���h|�k2`��;zc��`��6@p?_�!1�?� ���۵~o���d�֕݉��l�W��R�5�C�L\,�s���w��NRMu�U��=Nh�G#��'��m<5+ȧ� 1� �p�#5�xV�˿�s���d�"ݺ��ַ�{��Hx���je�Q��GDS�{1��Z1#�#5�|Xҿ��X⁝��n��5��}L^�F�Xܟ* ��������Òx,3����gs��?����Y�Vl�� W�]xt�[�r�9�a�]�F�ф��"q"�D|I�4�#ۍǌzWc{�4*�+�⹫�>]͵x*�l*�M��.E\Y��Ta}��nen1Wc�V��=iWkF�0Rz���L��*2?�'�R@1�t�kI���4�����w<_�1��]��V�1�������j�������Y����"�Rߦkt�0{��=H�/ތ�$b��mQ�R3|˓�c��@�G\�nNqߊn�܂=��� �����0?��/��B�� k��A!�~?z�.�����f�1cJ�r7~81Q��^zԇ�����%���x�B�ϧ֞�*�:�#������t�i����� �(�9<LP8\��6���sRl��\�����?ʀ�こH���)�7�p)m�i�����I���Z��T��c�K(��s��*0��A�k�� g��~;�� I���2˜� /ΑH�v�s��:T�����]�*2F{W3��l�V���ǵtv27t�JCF��sӜ��~\w�p� kB06�f�%^9��U��t5� {Ԩ}y�SD�#m��t�� ��Ͼ)x��C�/����5���^i�l�J!;������*6l��_\ۆg��ҩj5���!�ˌ�ǯ�V?���' �Uu��@�Ƿ�8�f�i�ݍd��?\�Jw��7�����ƫ�"��P*|�W�u�sܷy�����+���w�FÕ_\֬� ���oJʆ5����TN㎧��f���xsP�[��I����Z���&���a}BgV`1���q��ߴŸ�Yҁ�-ğ���?�� ��L������A�d~5���yW%ϼt�R�].v9*�9�Fju�.UpY�;�:X� �|d�o���q��3�ta#�)��?�kQ��ye����]�F~lc5B��y�sɬ��H���jp�72�J�B�S��'5�0�ٯIur��g;�?�=���Y��+༏!�q�ƾ��G}vR�1�V:���1RN�ӿ	<m�댾}̎;f�+R�/�� �`
�߀)�L3�7�X�<cnF+n�4���Kź��+(���<O��Y�?Z�R @��/~I��aq�x�QiZfj�5rg�l�e٤7lWc"Q�y�u~�� lX�?��zT�-jz���5���+ʵ��Z�2G��5�[�upGJ̓�is��zP���8���������+rM}��mq\���ě�w��#Uo�q�LRw-� �2O\W��l�Ew�~V��?�sT�G��DGi)=q_:|B����Ѻ�o"�|��v-��x5,h��ĸ_]�X�ޥ�r� ��1� }
g�9�E�#j��ƿhR<��]c?�~�~ɓ�Qnz~��%{T\�����T����8��p^� -f���V���j��ۭNˁ�1�:w�!̂���4��8#�d�N6�Տ�-r�G�̙��jFŗ�ל|db�\ex�#��iM��セ.����cg2��Y�Tx�����T��=p��|�����M�PN�m��+*s�.k����4���T
��W�rA?�U�݂��|�w7�-co�ҫ^|C���2ʯ9�8��fRrj��a�iWQ1��,)2�������4�է���֧�~,Xx����`}k�+�T�#`����d~��z���7a�P���?֦2��V��n}6�,�OQ�o�%�*��^?Ҹˈp���ڠd<n$j�����T�7�o� Z����Eld�~��j�z�VA�fm�;g�Kг���1�����Md��	�Ͷ4u������YAh��K��S�<�W�i3H��|�n���G1֩G����?�ֳ[�ãw��|X��N��U��l!�;hT�-�械���wO�G1ʖ�����=ܾ9�:Uk���e�?�����z�b������|��j� �$�vAv=+�Mu	��9S�וkM$vD�W�q]��fi4�=I�j����97sX����ͻJ����[ж9�`xg�6�r�����}+�;=�Q�;qR����c7J�XdUd�v���?�G��>��3!11�⼟⒖�v�r AV����
,����D/�� t��V3}�y��}��h�O݂3��#��F�Y5+�*B,ο�hC�E'�3�\nb�ϩ�����Pň��F��u$w�̰Hی��fX�O*����Kx�����{�9����_�c��+L��)�7 Nk�?ko�:w�;Q��a.68�}�s�z����:�?�v�n��x��'�C� / l�<������*��J&Q|�>$��~��=A'5����^���5k��� p �ۯ�^!����5�7w\y� ��W�'���zwß�æ���c&�2F2;rq�
�DU%gc⿆�  "�įZI6,t��ȼ������[>7�/��� K�'�dUU�
ۻ��K��Ox�@H-s'弜�Y��~%jW?𷵗[��o� )#h ?LM�8�w}��O�*xJ�O ū�˸gҸ�a$J ������ֽ��"O�(���3��0q�μ
�Ik��;�,�.��>�۠��zr��־���3kц<�F;�;�a�C"��mK >p�����.��E�Q���dg<�\s���g���A4�y�>]ͷ���r\�g�*�k�OE�?�l�V�%�I,�C�_Z����PӍ���O�j�ir�X��t���*F�3�@#5�\Y�&?��y��[��8UI�=<�K�;��+֬%��ۃ)PO ��i��IH�l����������3X6-#,���ن:`��赂�� �6vv�ef���Z`s��*HXd�g�].���r� �aX���'�I��o#�� �:�k8��!��j��| �c��d7lK?�:��i�KH\� �H�^Hw�޹��+�#b9J���f'��
�鄟/aHV3��Gv���oo,,nGR\g�kn��)#9 p�zV՞�l�`��~PzP=8ޣ'�֘1����*��#�/�݌v�E6�m�2��ݨGʒF t>�e����7v�ǫ[��O^���WVr���@�:�1���llV�w;��Բ��R��=j2���@,mg0u-�l�[��(�R�x��OJĻ,��v���hw�ʪ,y�P2��b�T��9ٓ�{�z^��c���ˠ�ȹZOo��P��{]��΀:/�;�y�����+������z�7�?��]w��G$�I�����Q���ԎG��:�9洎�r�����c�n�wOz`�
Xr*mQ��ѐ���Zlr#( ��ű����{�1}��+�o�g஛�7R����/!�w�RF0}s�
�jr��������	���mBḊ9�t��#��֐Wfu��_�I�^O�>8�[�6�`?v�T����{{׶���>�o�5ê@����D��6;��^��[I�~5����j���� I@��V����.h�����	�唑�Lw�����T��7dc����)���_�%"H.��3���  ��Oá�-��߉�F�aa�&�7���H�O��SR�L��짳��j����~c𯝿��wR]x�X���Q������G�R����\�&���	�?����v,Q����s4C�߽��� J�'��V���j�q�+�d3�����B�zz( }qYKFkt�	�U�n۰~5^dnpFq�z��������� �5�څ��;GZ�J��a��"�>Al�t3Z~:�}M*��q���U�b���4����M�8��1���$��ձ��p+�?g@�4��������0�6q�_q^��W�K��<���Yɷ�r�����.Î��WV/�m���#J�ǨX�<X1�n�Tc�*簮K���!��!�'����}�}kr� M޹>����/� �k���XɻV������5��� ?Je[�l2�k��l�#�@;S�
�wº=Mf� ���QL
�+���~�uYso�a��z������J&bC}�'�+�O������>����VY�1�Tg�>�k�?��������1C!L����4�����CG��>�'ֶ�a�-�L�U&�|�z�֔p���2����Ӝ�Ѱ ���x���5$����g�zr�~Y`A8�h蛣�Kg�������;�SPB��ܞ}jV��@8<�4}�� 蹏���c�L���~��m'�l8�_���N{9�<g�˖6p��bNZ��U�<��<��'��*���;�w���5�d�D6�(�� Verˎy�Y�Ԇ����W��7�Z &8�*Ke��}i��S�jH��	#+�@�?���X�7�	����\��W���f�A�s���~��Ҟ}gឲ�Ğh��_�V��&㍭����4wa2Ɍ4����4��F�����j��ǁޥ�@�~s��=:WY��]�R~��JO,ǒ�2q׭H�Gl㚻�;+���E g��������Ix�[��D�"�=����NI�����l�t�`�gں��sh˖�=s���:�6�y�7�<�_A�{Ė~'�"��%�'=A���wGe9).S��q���7�aִ��"���,��z�q�R9�$�O?�{��|M����I`&�Z�-
Pi�s�xG�*��+��|2C�	��⾉��<�l(l�\���Ԓ6CxU��Ϸ�������z)�3���R�ùb
�<u���ɗ�0G��8���
���^$H6X@߼?{'��ψ�0�� Y����J�n��}{R����wm�М񊨻�!�p���w���V��n���6�����5�`�V>�I���m�q�D��7�\�kS#X1�>c��#NI$���+vN�y�JV�����Y����y��Ӛ���s�Ե���O:h��@����v#�{g֓�B�q�ہR�m2g�88<R�����:� �@ni�M����9�"�Al��z����]�#�'=O���>^�2����I?�X������=}*��<8R/�(#�Jv�����pO� 뵆�� ]&����֗���Қr:�����.���=*11��68��GᓌsI���Ixi���|�dzץ� Y�2�:�}H<� ��y�0e(s���T�����:Ӊ|n��rFp=q��"��ݣ��N0|���Q��5�Z�+��Wm����#�� ׮��O�R`�X[oAҮC��Z�i��H�U���Y�O�*H�o^D>�	������Kɟ-qҼ��f�O v�^������@���O�9+�4��>m�F �����ɩ%��)�qZ"�P��������ў�\��R5�з�-�Ҙ�n�8�F��Q�#�k��+Ih�x-�@�,����^;�ݧ��5�j��ӱ��U�մ�*?1R6ܸ�"���p�w�;lr	��OS�on���M/��Q��l%�������6~8ӂ�p����9����[ݱ�v����8�zs�ۀ*���Ǵ@1�TM�O¶��Ԭ� sB�`ry��Yp��ڣ�*1|_7����>8�!M|o��}�iJ1W�� {
��"�V�<c <l3��A���q*�z~1ۅ���":)��B����ZU#{`p~����Q���h����:+x|���t����*��B��w�N�F2���R����z��~Rq�5��Y����%�>���Pѡ�џL��[�Ru�e�n����e��]�ۮ[�� � :ͭG��:��p1�jц�^:�kx�U�j[���=�t���0�WcB=��q�X���:P���+���v'5����p�9#��T��͵�����W�� ��܌�5��7��� ��t��jYH���o_(�)�&��$^O�W ��qRx�B��� ����4�s�sX���tt%�G��� $��	a��?�׹G���xW� ��Z�?�Z�UR	�Y�WR�M�T�T��j���@M9�?� �N�z�H�A�}*���v�W��]S&�����^�%F~��|L@�1��o#��*+Ī{���)�I� s���S�	�n��q]�~G�K�0Edf%����Q�h���˭66Y�g�+�*pQXQ�-�UZ�WoaUf_�ү����ҪȻ�8�t�}��8�R�m��wn��7�� �V�����4�Wnw)�q���cP�T�o��b�����o%�ڤu�$Q���U�^趰�ޣ*�Y�9�y���q�Qgm�?v��� O�A� 
�=N��9Վ�x�c�y�Wh�u�2g�ңa�y�[E)�]���}����kQӷ^�ԇ�1�Mx�-����ے^r0��^G����Ʌ;��ھ���
Iqk�%�=��~��5�kd
��s�=+CS�5-���Svã,@V����s^��ii��%����\W�[�MS���8р�=j�B<���Z���9�5S���CڢŘ~ �n��o��-� �5q�B��8��KVӚ�͐�����_.��>����D�"ϣ|6�t�n
lǞ�Md�|�K��� �l'��tGc�b<��v�F*%��jUR���*�#� w�^Y�B=��7c��T��}8�+��&�w=�C�@x/�3�|Fw��on�J�.O��^�\��'و��|~�M�w�6O�|#���Q�K''݉���!�ʢ� g�$��^{�ҭ;y���*���sڙ���U@�a�^����ş�SP�@X#l��9�ך󙜣+(�p�o�c�S^|8�V�;deT
=�==R�Rd��=���?��U��r�����Y � \Vg�M�W��Ōr���*��bT���F���۫]��f��q$g���~*�կ���V~!�f3Km"��˻nGZיlD"��zO�� c�5�W֒��6H�zu���� ��|I��^����!v(,� s�J�R��zm�V�(�����\��?l�kֲ��+D$]�aڿ�J\�l)FRw=C�N�io��ٴ�	���������_�^��|J�R�U��iK�0�ïLW��c�ڗ�u�58�$.řԏ�q�ϯA^�u�Mx���B
�}1�E%%ԮW�����6��{=:7Ve OO�"@������[~(�&����_N�>O.r�v��/le@9=k6�4��S��N��U�>8R�`7�.�:�ޘ�+�o�%��T;�ڙ�@d�֚ ��bY U��>��J���U7��q��ld�Wl!dP@$�<Q��6�y�v3�qү�RDхc��Ʋ6e�!�=������f�����s�/�l�R1��(�瞵B9D�K�GZ,!�j>g�qV��|��Xc�OZ��j��-��2m�0 �@����1��z�-��Ԍ�r�~���}��\����l�)g ��NM���������ң��F���� ���\Ӽ� [���R�������1�`S��f33ɝá�.�,���X�)�*=�[��[{2�?�5#0c�3L���%֛���ڬZHTp�9���Iy��=��]���B��Un.泾�� OO��Kk���<�8�Vn�-p�G=H�F�ɩN7��F��~in��]���ZRM��*w8�� ��̧#<��7h]A�rkJ��r�C��z�W&X4�UX� \�Ie0kq���ǽ���P �ֈ"�?����*��n�Q��UK]$<&G�ހ3f�K��A_b?J�K�c��2��ڶm��n���'�W�vĤ',���cc�`��GB}��M����T�n���x� �ul.mF�(/�/M��FT6r~�+������6O�9����e�;L�f���\��Iy��gYQ���y�j��L�?9�$ݨ9�2���`�����W��o�f��,�.�C.T�j��{��G���#==+��o�6~�s��{p����:��+���;a�p8#��~2�tH��h��+����R����� �͠�x��_N��`	)�}{����A�;���t��3)��X���ӓ�ҿ/�����$��p%��c���Z�ǋ��z�+k����#�)a�ӹ���sX��d��>|�t6�a6��"������fٯF�+o�kڍ�,�%�U<� 1_�~����R���� e<k�׿i�k���y��X�fa������B��G��v�I�U|@��� o.m^���)\�e���5���/�ҳ����� ��nf9=s���4 x��Q{��-2��#�JUܣ+���*�>��i�$cPQ��8�=��\�3�[�59#�4�",3ǵ���_P:U�;���H�%`��5T1�?LR�G��#�5�[�����f�"��U�U��^�%�S hJ�`�?�~|x_V������� ⾱�e�`����+c知sT\��w=D�"��-��5�ɮ���O���a����#ҡ���1�� ��\���!�K��q�iZ�m�H'5Ю����R���� �Wlt���\E����g���퉕��u��:����#���eԤA	�K��?||�|9n�iL�W����z�������u=R�K�I�U�1������bh�ʮ�?�w���K�KS��i5+̷�r��k��`7�BL[$���O�Ԛ��s�]4ϒ�����ZZ]��w��;Wl#�ӗ3��
�T0G�W�wt`�g�c�ҫ33>�EX1|�m� ��ϭhH���R:� +Bv�@O�jvY�<��E&C@0 ��e��q�#=qV,ˌ�9���VC�}��0?(��j�$}�� ��m|Gص�$~����ܶG~���?����[���3���迭}���� ��S�O�^|�gB'�-,�z(��V��ld�UXO�㚞i�?��(n՛#;1X�sޭI��OJdc���������6���ݙ�x��c�h�Ƥ� �s� ����(���_����2�u�#� � �~���KMcD��`J�)� �q_�,�Ƒ�]f�D��i9�ߥE��՗ہ֒%~R1�Ҳ���z~���p{�]�D�)1�߃��[�W$�ORq�4��P6O�ޕ����7z��P��{��x��)c��U��+q�r���@	�Fr@�Ȯ���,�H��UQڹ��6��JsI��#�(i=֎�h���tIt����G�lv%��j�ۚ�J��H~h���g���v)�=}�oagx�*��gܾ����"���q�G5���C�s��G$��?5Xmf#�=i���g��r2�j�VG4^�����<9���3]F������W�l$��Jۢ�ּP�&��`Ms!�݊��Fk����<�P��J]�ڶ�{�^�BrŎUKq�Uy$�N��� Π��!�zƤ�;x$�����*�����ԙ!���}�V;� �K���;u�T�̅�#ښ�������m>f1��)�'i�;�U�s�?�$��{�'ҕx#�''�x�y���@ߵ�8U��c��T���</a�)�F�}s����F�ڀ$[ƞA��犮�_l�_��?�*���i�n���/��;�7\7|�1H$v<Si�1����[֘o�~�0��=��Y�9�0N�>8F�{P>i�6���К���@�l\���ǰ9��יI*���'O�r �W����c��������"��境��dǜB�7�+��c�󞟭s����W��.O�WGk�Q��
BF���욷�j��*pOj�JϩD�~�$8=H8�z�]�N���z�'5B/�����7��t ��]�7�x�)���jN2r)� ᡵ��̿�'��>b����T3p�O[���>��]�7�Rh��9����p8���9#Pj/2����1O�ۜ�EB� ���4<��=�U���|������}��j<L���{U{?�Y�}�(�2����>pH�2*a,I�}R�đ��<��� ��
��i� h�F�I��	�ǭ'�lۆ��5\��DM�N:�T,N9'���4�A�R(����Z��E�e�G#d7pe(�*x�>�n����b�D��H�#��&��G���~h�eYF�/�횣p��޴M͚�dPE�*qhIQ*�ӵG=qn��T��+	����_�-�'��y.,��	�jG���ɦ�s�UO/�TP��>��jWVqô�G��d�$L����s�^���k}h�YA��Z�`c�U����Ռt qW�E��o֬)�Ut��VUQ� 8S�yߎ����z3G��W���O�	��K���>��v���*�9#ֽ�T�u�z^)�K�o��4!�|/�Ed�u�9ڳv�� \TV8Y�?7C���q�����d ~�a��rj�|���V�x�wȭ��d_S�o�>S� 
�1Ӑ����~��׉��6+c��@$?$� ���1�'�Y��\Ej}�-E�EN��@�V�:�/���9@ZU]�:�Zbf�m��������ln-rp]�|�q׵r�2!�Q��@�=DqM�֑v�ҴN����E+4�K,�t�;H͎K�O�W����s��Pq�MF�]��c� {w�l�b:
�1�� 1�j��F�F=?Jv�}(۾6Lg"�Â�4�p�=��	�6�ፅ�����I��]��t+V�,�8��J��qH��E��,���q�ߔ���P9=��i��pO\`Q` e�H��әz�Q.w}ܞ�Xsƞ_�����Y��W�#��^;a�@#��UX��ڣ�N�jj#oM�j_�jS�Gf��k���H���Y����ֳ'�3�b�GA&sRX�RT`c�U��s��x9�]#Y;1��'�v�.�Yr��s����n�SM�A�G�Ȯ�K����[�[Z]���ʤli{ށ���Ϣ��
֎�<>v�0``�+b<�;֑؎��TۇOʛOz��wd�ޕ���Qס�0����=�?�z���:��ˋw^�E4#�/�ŗÚ���c�¾���tH2ɏ���W�� Yc���O-������Y�O�����ZЈ�U �x�Lm�A�5a�=�
��$��43f2O4�4�ɞ��S��'�(�=I��D���zt��xT�	$�1 �J=S@���`3��x�FT2�RW9ni�w(�'�8��4A${�w%�GaQ���T��pO�����o݃���@�)��S]GA�qR}�=)���0)>���ۄ�3��~������LumY��̨�0�9�O���f\��H��� ��<�����a�ݺt���iX��\$���A�������}+à��4��cTڜ(�l���^��=r��Z��p����ֹ�7��1٩�����V�4�V�!\�v���^��8�sVE�g�����H�z]�Ƣ����A8��V�-E�!��mZ2A `c��m��t]��=h���ø�:���2�<���jk���*�i�c2�8��(ܐ���;�O =*=�ګ**��៘��]�X�`�TR[���A�@�ހ"��ʝr�3�Ү�A��ǘ��j�Q�2�5cT�j���P\C� �6��f���j[h<�ų���� g�'ˀ��9�����"��F��R��I�/'�鎟�M�iq[�-���H�B�mJz���$�l���Z���ܒ2O)/o��-G>£�>�?�!�ξ����N9�}?e��LFq��ڢ��c�Tqҳ���@��q��cRH�Fx���*��A
��Փj9�{格���S��@X��tlw��9Qbd��p� �H椹���!�"��0"�D�j�u�A��Jc��5�iV�2�/�/|A�|h�傻�Ҙ4k?�멯�VCl�x��Ӛ������w�x�M.)w��Y��8<g�_ҽ?��v��sod0��̑����?�u��U�\j2�L�[��� �V���2��Aw)�Տ4yaW��c�.p�w�_��WY��{v������_8���+6:dҚ�h��ѽ�j�r��^��ϱb��:6��P׵;8罺���P̪�� ���[�O�|9��%͕�� ���W���_4�� M:�u�f �����^��-SI�u���jkJC�E�q��>Rw6�3gR�I���=5�z]�E]��c�5��0��믄z�ݎ�o�C$���(?�{��_��$XG�xa�1���y���~j	��a`0x$�?�򤘮~T_Y�����|�"��+���۲�����Q������rf��9�9n~�ԡv��,��^�odb�s�Aڞ����:TjǿJw#��皠�n�S��ʙ y2��&rp@��"�*=)�|�XG�$r{��
�Wa`2(`qOX�|�����z��hmod��YW<�+���V�"�*�* Q�`W����; �84�h]OZ���-k��X�c���һ�/���VD�d�B�����ʾfk�1�w�|���C��5�*)��cQ�ꫯ�z�m�4m����/�:�PR&�v_@q^�/.៘�����3y�0<i*+�^�]��� �u-��B�#i�OָY���.|ۆg��<�3W���6��}9=}*彺B䁂:涌��Rr܂�K�F�?
�*�ۢ(V*0J���#=ls��1��${�2�3�X�9�I�F�*Qۨ�KI�u��H���H���O+�v3����@�g���i��#��ǵ?v����8�h4;z�=3�V[	f����*����^G
��<v�mj�)j>� ?�����N��k=s;����<� _ֿBt�<�?p�pp?�~|����X���Y�`��c=V���Efr6��Ҽ��l궃���߻z�T�l{ՙ�ç�X�؝��"�_�ޥHˀq��q�R 㷽 e�M,J[�&��*�Mh@ �'�>b��9!�\g#���^�;o
�@�գVZ�Wn:6�� *�'��=�x����/����������9�k9>V�k%t~c���C�����}A� =iż�F$��w�N�tۍU�N��˖��e�H�R���P?��A��U�A�)�Aێ=i͕P3�d��#`F2�:��������ژ�0i�����J�`1�)?z����ӧ4�F�[��<�\Fv����7d��ND{X���e�c�����Vݕ��j\�.q�9�H��c��0"h����\ӷ�ݤ���N�Y�d~�v���"��ӂA��3C�#֍�1�z^:c� F]�s�Rn
�tއ��=:Ӱ ��Ҁ���֗y����4�9#Ӟ:�Cn��G�?�r�e�'n2Tq��)��n������fX�^��?����4Ƭs^QQՁ����nYK���. ���N�������M=�ƨ�zg>�S�DN�S��u����:�JQ[�������zY$��l��]pO�=����zU��8��=� �\�p�)nON��`#8�~l�S� է={Sʃ�8�J����_J@7�X����# sR4~Y���j��e$g�4 ��X8�\t�R����l�X�Uvs���K����N�+�U�2A�N�[�D�m�pW�A�y�O�����^��%�_X���;�	�L���M��}%1ci�Bm� �y���~R�s�*�ӬC�����j�m���EH��-ץ\�ET�<
��f�Аw�J|c���:c�r���\o� ��g�@�g���G� � s\ּwH3��nA����K�,D���}@���s�Rx�A�v���vȰ>Qx�N~��~�x�hS�3��׵~O�d�/ōqqʿ� g�E9=P$�sФ��|e����G�1��PM�\x�A�\8���d^A ����b0qG3����j��� ��.2��~����^.XĎ͜�FH�^My]Ϟ{|�Pj�M�	��q� �v
ǩ���ƛ[�"E �@�=����_�$ۛ�$�߸��^6�6gv��~V8�F�hz���g�����9��c�~�ߵ7�����3�bBA�b��ƪ>\>�� Z��<v�
��~�6��>�>p~��M�I��N�����M77s�=���F
���='�Gƹ�j���!���Z�ߴ���� j��O?��>�p۰;�d��~���|~��5g>�\�?:�O��1�s��n��?�p�"��W�Sʆ`ű��Q�;���p��Qf^C|���u>��|Ak�&�y<�k�7(�)����a�u�9��堮}⏏����,དྷ0�����o�_`�7���d��|�wz�� ?�~k�)M׉����Q�����_ ڛ[=.:Fc���\��B���\.s��Z����_���,7S��� \V�*c��U�̷�Ǌ����V�@<j03� %�^4��9AɯER+�<j��H/a�8�E� ј���C�C&pkԵQ�۲�����n�0
O=�)������~6�ڿ'�ǁیW{���(<,#;Y3�#���>$)������ �1T�q��0�~8�����:\�T���3�7��>���׶C��ĿdIC�'�v�������%�d��z���jT����C
���*�IӜ�MY��K�=��~p{S5"��;W#�k�,-^��D��=��u�6#�5�!3�N��F�zt�����6�㗄�fhd��6�p@�< �� ��M�?�~cx�R�_j���X��Lmb	�_��׳�aD��c�4]��ӿ�_>�:�j=sT����ZC�J<����%��ʭ%�@�U��u+���7ڙq�O�4�����q�������X  @8�Q���f8����V�?Z��mB��RiGc�ң�e�)&�ᇻZz�ʏՖ���5�h���O�~О�6����Z���m�#2�B�(���+j7���.}p��i]��?R����Z�ͪC�-Q��3��	]F^����ۮK�����ZU��9���3�d�zR�+��D?�G���}@� �O�y��HC�5���˂wK���F��ATku3��ه�i݋��������/���ˑ�Ȫ��LxCi��A8�>�2V�}�We�M��M���2Jwuc#?3M��w���H?�c����R�S�R0O�*��N?.����k1b�0Q��J��$�)���?Jʏ����*�
ϼg� >�8�>?�S¬��$8<q_��+�X���Oj�%��Vga�Ecד�~��d~�'�%��0�(-�C.Hӥt:|�q�vC���� *���X�OY�nXL���џ[� ħKSˈ�$��Eq��Ɛ���A�g���ڋ���F�T��U�m�ZGb娇LՍ�V�N������\��G2�^G�^c�+�=dc���&�BO��ω�4�6?CM���x��#:�=�=~��K��l�x��}��YB�OSl}�\��� J�:��G��٭�I#6���j?��_^�/ߓ��QڂlC����
 a�z�Oo��w��Ny47��@=�I�7�9#��9��2p=�g׎���I!�@�Zd�����T3�}q�����W_g���xǥ@��s/@+cH���f�?(����I�b0L�9�dpO������֢��c����1�@�W<��+N:ݰͻ�Y�O�M��Up��Kq��b�����6��_g�ͺž��$[��$�?Ŏk����q�?^���e�T��~�Ή��bC����?I$�6�p���*݁&�iW�m�3�s���5��� 5���u#��"���0�٨���b��_-�߼A����)I�3x����A�Uq��{t�[������4�7n�X�$�u�K�:�'������(>�>v���֧��>����d��[�bެ+Z�]Ѯ4ϖ�!��*���5�o��K�xN����^菻�5��s\;�\;'8�'�Ƕ1U�}�s�v��:,
��#}Z�i�9Тfs��n+�%�&k���Q���/�,�Y���������?P��7��,n���� ԷZ׆v��U}�?�~Z��mr.EԄ7=j9>+kXa<��O�y���Iw?Rc�<=�[�DѪ�-��֨�k�L*\\�G$�䯵x��������V��5��r�z�}+H�Z���h�26����8+����]�]�G�լ�P�	���WW2=Fj�Z���b/��ٜ푎3�?G�]��:>6�[�+ö�I@*�ne@�z�:�99~տ�z����ㇳ�;^x��l�����O1�����d9����nj��6����-�{O�k������8�K�ۜ�s��W����  �HcG��}�˹�W�<5&3q9뻥]o�f8ԉ�-��[��ď����~���N�P��W�O9'8�'N�R]Y�8�>��\�Q��������9q��?L�3�%�hz������`nTO��K��ݚK]���R!X��F���M�q!0�l��_R֬�9��jvSXC;�*� ������G�����c�W	i�	<ֳ�V���q���{��^{� 6��4/��C�w��I�I�ξ��T_R9�#�q	�k�=1>'xy�lw?�¾B��<m���1�
y�׆Y��V�C��1�j���]kK%ԥϣ��ԩ���r���}�O6�q�N?,�]�Q*E�L
�[��� �)����ֺE��W<�x�4��\�Ҝ0��&����?\��7��<�c�ޅ#�������;q�,�4�4u��FU�=Z��W�� f��2:o�YS�s��D�s�$c!j\S�U�sq~%x���F�h��s��Z����j����$񁀬0:c�k=�����돥*�~�4�s3>٥�bd�'��1�#�$P�})�n�c�ެCv��3RC�����9�*� ���g��*�o�t88�H6�g��zP���^����2�p=(��[ �3ڣ�Nr2W�Zk1�NN9�o����8�	Z3���zTO�rAb���S�Y �In�5��3� >� 6}{ӕ���$��{a��zT�f�r:���PE̒|��{��8��̹uj��q��*��W���F��8C��矧��,(YYCq��v�X��_n�{�FF�q����i��8(�?����}��ӑO���#�v�qMo��8ȥ2"���s�@V�y�F�b>nG���3�Cu����9�s@�6��{w��翮A��5�Z���㷱�㕮+HI sɢ��� jb�b���y���U�x·�eo�g�p��m͎�C�f\�6�n�mcF�[�#0�$����}����ڇ����*�m�	��1n�s������
�K#zq=����#�_�aSIz�7�3��+�U�HB����`ґ۠�:STrN8��,�P���&��Zu�"��y�m�����fȌ�%ۜ�b/o�x8ǽ@�	I�JU��$�(���Ja�f�.A&�gˌ�>�7��R����a��n���Qm�7�a�s��.A�c_4��њ���� ����ї~xG�?xL�|��d�X`��}޼/οau=�Q��	������������&�x�΁3��P850��vd�	���+hV�=��z�A���\�-s-���4S�
P�z:����g��k�jsXb��-���z6O^��UY��z�Z#T�H$�9�"0���l{��m`ŀ*���8瞵#)���aSD��N}h�+tě>Q��í*�P$��*]IV��f�;TR�#�����_֝���F˂A�<��A���q��eI��K��c�c��5 D>�n���V��Tݥ6��é�ƞi� =7q�0��ă���Nh�RF��q�3q��˝�#�>��V8`��=9�#v�Y@�N�����8��qV<� ���횁�n�:�M $lw����22*fSp�S��y��H���3���Ҥh<���� *��1�?1����3.1�c�Z3]D,c�g̜��Z�X2�t8�M  U'<`7a֝��2��v�ӟ�J��O#�GRO�y�j��$�-���aP��S49n?*b \�?�h��9�T0s�)�[�,3�c?˥5Pd�y�@��4h2��*3��`�)��8�����R
)'�޿���dV+2,y��Ұ��eH�>��@��}v���6��	C��ND;���$��1=�[ߊ���_Y�೅��?��С�pr9�� �le�uds�g�3�� 8��ks��C;��#� L����Z���zn�G�]�?����� ?�t�/+�z��TQ�l
� �5b3��}j�k��y�YR�Hg���!m��U#i��э�BG?\W1����v�t������k.���֑ �`?�O)#8\~��M��1k�Z 
�NCd�oֿU|gj�$�fUےNF:W�� �1z�|WԚ�E�A��	��ߥ)n8�q�"�ѕ,p�Ճ�HFK���ׂI�h��l�����Y�0�g�I�,�9 ��j�u��.On)�e]�X����0+�����x�s��+t�*��2:����`�n'�)�63�?W�~�z��x�9���c����D7cʗB�䍤�����3��gZ�����G��~�i>�C��xz�;{�8RU2��z�¼?���e��9����f���H��_�z�G�5|����ך��۵��3���~?Z�Mҵ-Z{[9.%�)���?����߳�ֿ�w_�y����^x�W��¾�<M��F[�H�mŁۜ�q�t�_ʫ�N���bXnl�W��[08+"�QD�n��0��s^��bkz<�$��+u�==�H���c�5������
�Me+#D�Պ�>V$�>�t�w(%��1��E�A ��>8�(��6�֠gG��ʛŶh2x��G�?:�B���M1� ���}F:������t�9�@���R��`�#�� A_�^�����S�<��ӎ�Ұ��7L��~����k[)T�O�YG�\�q[�t��О���#=*U?)��ڡC���w`�@G�I�=񔛮��Е��1ڼ�Ő�zO�~���/T��9�p$�6r��ק]Z��Q�a^�E��ɕ�5�~��:SB����9D������,?�Y0ܙ�X7��� �µ~'j�w�u�l��C9@��'��Er�HY�	�0�j�Ʒ?V�c�7|/q��r?�^�o�b�ׁ~�Q��*��zd~j9�~��b@�8�%u/E�zb�^�����c�U���v챦n>` ҷ�MR��T�5a�S��o�_>�x1� ,�?#]�|��5��P_����� ֈKs�Ōc�7nv�1��Vt�]�Q��hx�E���Tt�c�l��b5�I�j�-�v&fP���j2$Pw
���h��/ Vm��h�3�)�B����?�7�s�g<�g�Ӧ�F�����f�9�N?>	��v���]�<1�x���m$�`>fT$v� ϕHR[�z�o�o���τ���U�Iz����#��=(V"M��վ��H�3M�\��,�Y�VO��/�x�����Y%�C�E���z��#�E����si1[���ʓ�W��:����e��ym#��巪�?(a����AZr�=��򟊼��6�(�K9-��*�����>x��MK����&]�V2F:�=+�_��\��<]��Y۬o$�Z�
NG8�+��x�N�G��uY-�Y!�b����>��_3I>�愖�u��]F�J�C�Fs��\_�=�Ծ-�}{�z��Ț�/����1Py$�,r}j-[K1�8�FkV-+�5rHOrI��EF�R��oʽi6���̆;x�F)�[,s4A��8�)���"��;����{wYK�_�Z �|�|_��B�+���Q�vv;Fp8�<c�W�����x�Oے�!��s������[�x�ic#�. >��\�~#x�zޘ���� �hN sYH?gNkf ����e��Ts�Z�.��E��c�4�ķz�Ƽ�₏��8�?��No��f������:n����@���|/���~��>د���^A��� 1� W�� ����z���O�t���Z� g�^@�D�+~����ϡ�y�)�N���S�z)���M��������� ��	\���Lo��Js)^�i1�`|�֝��'9<SX����v��M�2Wp?�!��,���`�S �'�j�)��zP�wq��� �cy9�⑔g9 S���z|И��@�Լt��:�=)�9�G��'����rhPlS�<�L�b�(>�u��c��Ux�V��k^O�Wo�Wo����1E���#�{S�]���/ �ֻ��j�kr�6�1� Ҽ�KUa���c5�|r);pGOZ��wb߉�m{⋦�����U��������TR���δ��yd��D��&��E��3Q�+#�;B���{��r84�&G8�ҁ�^m���su?�T�-� �>E*�<��ۂ:� ��;���{u!�m`z`W_q�N�wpҸ�3NO�xg�Ą����tTuɬ�"?S��}�\x�_�L��&hb�|�]Xe��F1�z��K7�V�B]��.Ó��\�OHq�?�z���s�>�����Ǖ��7p�p��9�Tc����r0�3�V���|�+�sU���I�s��\\���t�?N��ޤ���_
��q�3һ�j[ōJ|Σ�!�Z��\�8�P5�_0ۏL��Es��/ڿ�Z֟%������W�ּ��'V�{�ɤ��F��+n��=J�����1�ެZ��d���E!������FGV#=2*^d��mQ�N?:�C����h_a�xP�#�q�M�q�k.�4��zR� QI�c��`P7Ϟ���)&��B�͎��~�ʚ[3� ��M����c4�-� ��Dp��kh�����p ���?�y�\]ȿ,�v��{{P2����g�Un}sCq��i�>� w�?�ӱޅ�Q�u� 3Ҝ9�8�$P}�#����@�3ޚN}�F�����r�b���F� ��&�����I3�RA%�s֛/�9�jkY�J=W�>����Dֺm�6���:n}c�TLg��J��A��s��)�B��)p��zt�K� ��@UUbs�>��f�d����?��S#O� ~��{đ��Z`Ap����������@�3�1�󊍀Rz��S#|ˑ�=?�J ��������R}�������fTBU[���>�^ǩ���q�@/6���ޚ�d��Jo�=3��Mq0nT�J �V� X�:�����(l`��ۻ�
�NO�ƴ�M��S�QT*{Q�!��Q��|u��ܚ��-|?2�Aw�0�h� ����c��n��MJ��kjW�j�k��=;��������?�Z[�nDѧފ��A ��_�����1�d�ƿ�d�4��@�:��u����=׮�� k�o������L*t���h��*.�`:Sv���w4 �JG^�2��v���#�0�.>����E9�A+n�1c�B�Z�zUЪ��z �����j6]ŏ�y<p쐹?U)�>�`� ^��[�<R�I���
:s��[U7�(����c���&p�`g֡��r8�ǵ��d��QO�z�n���5+Ya��e�A�Vb����~�������ng��?d�?4��4k�ª��?�O��o��M�j�}1'��~�4�p��r�.�a���7K�h�ʑ�^})��BiH����[1�@<�o���s��Z�_��[��4�:d��V� Î?:�?~��!Фc�o�F]G�ZF�s'ǔ*g'��c�#�jӻ�n����O��!�G�P���Ebb�����&?"k^e�\�c����^�p�4�$��#3G;<h7`����6�T�̓O4c�oU��E˸r2/v�1AO-FM=�X�|�ȧةΞ�q"�"o�';��֗2fȼ���=�;SV=���ñ���F�%FB6��=�4,���J�ǂd��d9�����0P��������ۄc��z�j���I�`a��/��T-
X�`8'�9���ݫ~K�� QR4������I��Kkcqt���d8��@�;�>�q�n�ȸ�h�A��D�$�}i�N��j?��ؘ3ƨ�|JU���v"8����ߚ\�\�?;w�?ʜc���n1N���h������Ӗ��N�K�S���9��\D�����y#�+��:T�J�nhd�B�*si7�9	���s�\˸r2��)���03�jn�3�HW?��9�`Tz��M}*�<��?ژ���q�6A��$���}i�8�F>l��Z����"dۆ�o9G����&�X-�Wz�׿�G�A�T�ƪ���z�w_ץ9����H<�~�DԔ��v������&�ͥ�HĄ\}���gӡ�λ���v���9�?Ɵ��� ���)q�n2�����S�����)s"�Pdn#��'�k�>����D���~�5�aj8��Bq� =G�_�|?�Ho��VH�~�FJ9�
�q�� ﴋ�Щ� t������x�}k����mt�!u܍`�;s�jя��ӗt��z�_銞ep�gұgh�N�e�k������كi7@(����M�k�3�4�u266���̃��Vnl�]�nH���A���?��30U����$���u��H��/-t����N@�`1�Q�jyƩ��fA̋��J������� ��_Z],W+�_(����?���v�r8}��Z�g����|\_#R`-�s�`�_��U�.Ti�g�?j�x���{�b�F�ݺǨ�&�k�J�y��3\��i�:V����`�	:�~�sG�"z�(e���% ~T)���u��I�⣑[q#�]~է�b�v?�� I>�J�DQ+�v֐t�꽠��9����q� ֧6N}z�޶����KXH#��9�i#�.�6ұ&3���9�̃ٳc�A��Ӽ�C�ku��Fq�x�zy�p~���A��~V!��|�^���ݿ�r=�k�>�<U�3&YN '�[����p�cX�-�:��:~��_�w,(��� $���UFq3�d��1��ºφ~-Y���ʗq�FW���}+�L�X�>��5����~�� :���k��K��@�#^kǴ8A�ݺ�3��|��3�ڟů��n����o�X8B�+3|�%�x��Z�Ek\ÖNW=�� ����3��
r9�+����x�]yrDL�.�����z��/�E��i4+M&Y#���
�T.S��W�~�z�t}F;�7��a'�nW���Rmw����2_��(wV�=��FN�\�ۍ� 0?
���O��^0��I�a���3��~l�k�c�k��Ej����˙J���xFnH#�d��3ӏ�]i�Q�(��������>�b��(�v���.Z�t�1<xt���>W���<W�¿h�%����y�R�����'������$�Ðq�8���^2���C*�Q��Q(�#�튉I2��[%FE��1�+V*>7
��� io��A�ۤq�$�᳁���+�����̄Eo
�8Y�N���X�g# >���������'��%Y��U�ؙ8��j6���%·�Āq����]��康�O��x�T��w�O<h�3�� +�I?h�
�3���_ָ���_�?Ȓ�"H8q�ҕ��˹�'į���^�X-%7wY�X��j���W��O]\F�ղ�"`A�nݫ�~/�q%��$��~�q��֙� 
?�С"uP	�%^~3V�pp����������R۩��60p����5�G�?��wkt�o1፿֧��'�8�@����PEȕ��?O/�<d��f$�� ��v�;���e[{���ٮ�
�)��⽶�R���Tlg�ڎBF֥�ʳ#�!� CV��
� �¤�V\��o��Q�֢X����� �!iH?(��&��m�yg�q��o�+�P�'�7���Dllr ���W��t�v0k�O���z�������h�9�y���Ҏm4c���~�xu�{Q��*.�`�v���=�������� �̾&�}�\EO!]px��~��*e.!��3���h\���j�[$t��J�#"�^K�M{����Y���#��~�*�ɾ*��'��T� J~ЎTx�%��0:�RB�����+ؗ�G�Z��{o�L�0O��H��� ��;�S��S�^p8��)�wQI\1�d��~�y�/	\j�N~�}�(,p;�k�_��Ѩu���d\f�K࿀�Q��	ݔ��ʣo<��j��=I�]���$�^�������Apf�N���=3��ZG}{��{�`��h�=BW���&�ki�h:e���$3���,�[��x���(������>y@yϱ����a����ߚM�����u����W��W�~��%�~�z��2$A�
�1�/j�><xWſ�=>I���KV%dYGϟQ�v�D�ι��;�ƶ������}�~n�J=����R��g�_%�"e�������y6�$�w��y�?d���R��>�o\9-$L�N�����c��B���Q��k>s~S���݆�p1@�u�����{��1��c�j�۶��RIʅ��|P�O����鵺�΃��o0n��y�Es���z� �1�Cg�=E���-�3`-����� ��Ή�<��2m�f��� �`�u�1���_���=6A��^��񯉴��+ĺF��B�pۇ�GQ�W�o�A����}�F�x�\c�z枬���FV�0x8���ˑۊ���v���ҮǭD�`�Ui�fl�'#��.Ӵ�k4k�/\�T�עs���\³/��!��kʾ'@Ӷ���
�c�G����i��6��h*[q֟7a�x?čr������3&0��O
�������޹����Pz8�+�_�����~#^f�TE����c��� J�!��u�P�T���2�N8��w���Fۏ\t�LGS�k�v��uu#�a�ʉ��Q��M�u�����������'���0�;�Zll���⾢� ��.�����ď��������C�Ŀ�;c�ү�٣�I$\�n�rx���U��ޯ�a���i�������� ���2�^,�]��� ���F�2$���Hz摤^:{d~F��� ��nV���|�� ��0�º�"��m�䴹�ʏ�� 9��j/3h��G�G����Ō��)���)�u4��^1��v� 
|�ʏ�r��{b�_$�{`WԿ������\�wO�B�Zg�0�������2?�>q{3��pF��T�ȫ����_�N�iΫLs�����4�������L�l~X��>T|��l1�ܑ֔�q�����K�_�+�w�?�/�0e�`�Dǹ�O�B*����>Q�+���U�o{c�}h��lѨa��y� ����P��M�������� ��^�$�������'i��pM}f`�@��r0~`�/�0ˍڪ��_z^ԮT|�!�A�;mδ�P4!�'�v��W���"��8r	�kž2|'��Ž��dI�9Ƕ~�Թ�q�y������~cڬB�'����U
���
�	��b��i���RnqP�&�
�|�p g��EKqbo���#����~��� A_G�/��� �?�a�.�m ݕ=8��v��ɶ=A]A�3��Ys�(��ȑɑ��S��d����� �g�CjA��8��#�����yc��:��>r��)dU�q��������}t��y�f��yo1���z������?�W�0$�֏h/f�� �np�SH�<̕#�J��o�'���U3�G�ӓ�	�#��&Q8۟qG8��>CBd�cBI�pH�h�7���3_a/�<i��FP�~��V����@4s�*>=Y6�r6 �\sG����f��־�_�'������)5j?�'� ��X�睪G����,���߅J�*.I c����-��qHĶ����n8�s��O�'�-!۪(l����S��^�w>B���?�4�v�d��?����;�W�2����o��L߰RI���9��r�@����*>9�M��8�S���%H��J�� ���ͨ¼�r�!?�R���ЮN����,���0�G�_h^C��^��]Ƹ����O�0*]J4��I��o���P��RG'�Z=�T|f���"���*�3lc�@Q��W�_��6rG��q���0� �sI�k�F��h��\����V$��|÷*	��k�����x��(�΄��%��	i$b6��-�e�<Q�r��� ;kc�0i�q�@cǽ}�� mԠ���*��Ѱ��:����ч�]ύc�N�w��?:o���r��������	�ot�>�0GO:B?*���e�� ��S�����i{F�w>'�`��Nx-��i�y��.3�1���-� �Uu�oL�� 2sT�� �|�4�j�{��ߙ��f��)]�($z�i�MjT$��Z�i��v/�j���G�?��v�p5�����~��^�|����)�3׎����I0s��+�?���{W�7���͟�s��e� �}Zn*��F��+ (��ʏ��.<���,q��O�f��<����?�O�E`TQ�8��V#� �{i�>}E=Է����_$|Ի�lA#wu�� ���� �x�?x�c� q� |梓�	�1%u���?��?h�Đ�vYXg���F�	�Y��q�5��?�O}_� s��'��^��	� ��6�o�z�_�K��Au>�#�����c�j�W6��|��2B+0��~��?�_�m�>sy����?\פx/�G��� �l��C�T{Ar�l~lxW�>)��6��yy4�t�2}Yy���� �=|K�[�/�a�.�j��xv����"�����t_��N�����s۵um*��  � `
��ȣϾ|��>=M��E\=���H}Y�נ_7A����>�d�ԣ2ԕ����
�o��#������l�^(���u=�胫�A
���ڧ-� zf�j�� �ӛ����*?��,~f3�}(�rTc9֏�m�1V��Hn<�I*��j+��u32����EXa2d�Z�} X�Ȩ�U����֡���h(��PK   [�Tqn�D       jsons/user_defined.json���n�0�_q��0`�k����vӲ���jr�t�R������Lӄt��&�E�����s��d���S������$�'��e�x๞�'U�l_������?���;'�d�7��u���E;�:e�g����1��b�^(��fbx�$qF��CB�0]�i�y�(�ss���p7tZ���4#U�iYo'���M5��_�W��ș=}���~F�r��gl%m������kݳ��}"!�����nQS�ߍ�Bq��kN��v/�XEۙ^�U�
<����$���/��N��'�b�n�+�$���7�~y �{����:п��)� �1 XJ@ bc�	�P s@�ԇ�~d�+�#Y��#�>:��G� u �3� J@2tF���e���>A� ����B5����Tz�G"5���"Aw����cf`�B��=c�P>��c�PE ��_y���vF������#c������1`�&�V���K�/;92��d8b	�T��NF��(�VNF,A]7}�ɇ�B��֗�|���$�=���0��;@�	8��;5���{;�5A6t�K�f�ܤ���)��2��&`���v�vHW��W�w t�W���k64՟��.?�=~�/!�]��*���%���o�>��7����/�F�#�₿qV^��C�+HYax�o'��Uq���ί.��IZ3�ӡ�i��I� �9�@�Bi���HѡБ��P 7y�s�A]Ñ�]v�؅}Q}ݠX��6hQ�����A�"4�_��A��D�<1hQ��>;k�W�ls��5VΡ�Q_��L�Ư�3�����n�PK
   [�T;m7�  ��                   cirkitFile.jsonPK
   *V�TD�98- Cz /             �  images/ac84e508-e9ae-4a97-a513-a57c89513e93.jpgPK
   T�T_��jOw  � /             g images/cbe86463-f5ee-4cb1-a8cd-cff047d8f75f.jpgPK
   [�Tqn�D                 � jsons/user_defined.jsonPK      <  |�   